////////////////////////////////////////////////////////////////////////////////////
//Module name: Top Level Module
//File name: simd_top_level.h
//Descreption: Top level module for SIMD unit
////////////////////////////////////////////////////////////////////////////////////
module simd_top_level(
	clk,
	reset,
	valid_data,
	valid_instruction,
	data_size,
	data,
	valid_output,
	out
);

	//instansiate core control

	//instancisate MC

	//instanctate Memory

	//instanciate proccessing units 

endmodule // simd_top_level