////////////////////////////////////////////////////////////////////////////////////
//Module name: Top Level Module
//File name: simd_top_level.h
//Descreption: Top level module for SIMD unit
////////////////////////////////////////////////////////////////////////////////////
module simd_top_level(

);

endmodule // simd_top_level