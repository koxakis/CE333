module alu(
    clk,
    inA,
    inB,
    opcode,
    result,
    extra_result,
    zero
    );
    
    parameter ADD = 3'b000; //0
    parameter SUB = 3'b001; //1
    parameter OR  = 3'b010; //2
    parameter AND = 3'b011; //3
    parameter NOT = 3'b100; //4
    parameter MUL = 3'b101; //5
    parameter SLL = 3'b110; //6
    parameter SLR = 3'b111; //7
    
    input                      clk;
    input       [31:0]         inA, inB;
    input       [2:0]          opcode;
    output reg  [31:0]         result, extra_result;
    output reg                 zero;
    
    reg [63:0]     total_result;
    wire[63:0]     mul_res;
    
    multiplier mu0(inA, inB, mul_res);
    
    always@(posedge clk)
    begin
    
        total_result = 64'b0;
    
        case(opcode)
        
                ADD:
                begin
                    total_result = inA + inB;
                end
                
                SUB:
                begin
                    total_result = inA - inB;
                end
                
                OR:
                begin
                    total_result = inA | inB;
                end
                
                AND:
                begin
                    total_result = inA & inB;
                end
                
                NOT:
                begin
                    total_result = ~ inA;
                end
                
                MUL:
                begin
                    total_result = mul_res;
                end
                
                SLL:
                begin
                    total_result = inA << inB[4:0];
                end 
                
                SLR:
                begin
                    total_result = inA >> inB[4:0];
                end
                
            
        endcase
        
        
        if( total_result == 0)    zero = 1'b1;
        else                      zero = 1'b0;
        
        result       <= total_result[ 31:0];
        extra_result <= total_result[63:32];
            
        
    end
endmodule

module test_alu;

    parameter ADD = 3'b000; //0
    parameter SUB = 3'b001; //1 
    parameter OR  = 3'b010; //2
    parameter AND = 3'b011; //3
    parameter NOT = 3'b100; //4
    parameter MUL = 3'b101; //5
    parameter SLL = 3'b110; //6
    parameter SLR = 3'b111; //7
    
    reg[31:0] inA, inB, out, out_mul;
    reg [2:0] opcode;
    
    wire [31:0] res, extra_res;
    wire zero;
    
    reg clk;
    
    alu alu0(clk, inA, inB, opcode, res, extra_res); 
    
    always #10 clk = ~clk;
    
    initial
    begin
        clk = 1;
        
        //ADDITIONS
        #20 
        inA = 32'b11111111111111111111111111111111;
        inB = 20;
        opcode = ADD;
        
        #20 
        inA = 1256;
        inB = 1453;
        opcode = ADD;
        
        #20 
        inA = 2018;
        inB = 1997;
        opcode = ADD;
        
        #20 
        inA = -8964;
        inB = 78965;
        opcode = ADD;
        
        #20 
        inA = 0;
        inB = 21230;
        opcode = ADD;
        
        //SUBSTRACTIONS
        #20 
        inA = 10;
        inB = 20;
        opcode = SUB;
        
        #20 
        inA = 1256;
        inB = 1453;
        opcode = SUB;
        
        #20 
        inA = 2018;
        inB = 1997;
        opcode = SUB;
        
        #20 
        inA = -8964;
        inB = 78965;
        opcode = SUB;
        
        #20 
        inA = 0;
        inB = 21230;
        opcode = SUB;
        
        //OR
        #20 
        inA = 10;
        inB = 20;
        opcode = OR;
        
        #20 
        inA = 1256;
        inB = 1453;
        opcode = OR;
        
        #20 
        inA = 2018;
        inB = 1997;
        opcode = OR;
        
        #20 
        inA = -1;
        inB = 78965;
        opcode = OR;
        
        #20 
        inA = 0;
        inB = 21230;
        opcode = OR;
        
        //AND
        #20 
        inA = 10;
        inB = 20;
        opcode = AND;
        
        #20 
        inA = 1256;
        inB = 1453;
        opcode = AND;
        
        #20 
        inA = 2018;
        inB = 1997;
        opcode = AND;
        
        #20 
        inA = -1;
        inB = 78965;
        opcode = AND;
        
        #20 
        inA = 0;
        inB = 21230;
        opcode = AND;
        
        //NOT
        #20 
        inA = 10;
        opcode = NOT;
        
        #20 
        inA = 12354;
        opcode = NOT;
        
        #20 
        inA = 1997;
        opcode = NOT;
        
        #20 
        inA = 1994;
        opcode = NOT;
        
        #20 
        inA = 148952;
        opcode = NOT;
        
        //MULTIPLICATIONS
        #20 
        inA = 10;
        inB = 20;
        opcode = MUL;
        
        #20 
        inA = 1256;
        inB = 1453;
        opcode = MUL;
        
        #20 
        inA = 2018;
        inB = 1997;
        opcode = MUL;
        
        #20 
        inA = -8964;
        inB = 78965;
        opcode = MUL;
        
        #20 
        inA = 0;
        inB = 21230;
        opcode = MUL;
        
        //SHIFT LEFT
        #20 
        inA = 10;
        inB = 20;
        opcode = SLL;
        
        #20 
        inA = 1256;
        inB = 32;
        opcode = SLL;
        
        #20 
        inA = 2018;
        inB = 14;
        opcode = SLL;
        
        #20 
        inA = -8964;
        inB = 556;
        opcode = SLL;
        
        #20 
        inA = 0;
        inB = 21230;
        opcode = SLL;
        
        //SHIFT RIGHT
        #20 
        inA = 10;
        inB = 20;
        opcode = SLR;
        
        #20 
        inA = 1256;
        inB = 32;
        opcode = SLR;
        
        #20 
        inA = 2018;
        inB = 14;
        opcode = SLR;
        
        #20 
        inA = -8964;
        inB = 556;
        opcode = SLR;
        
        #20 
        inA = 0;
        inB = 21230;
        opcode = SLR;
        
        
    end
    
endmodule

module HA (I1, I2, sum, carry);
input I1, I2;
output sum, carry;
xor (sum, I1, I2);
and (carry, I1, I2);
endmodule

module FA (I1, I2, I3, sum, carry);
input I1, I2, I3;
output sum, carry;
xor (xout, I1, I2);
xor (sum, xout, I3);
and (o1, I1, I2);
and (o2, xout, I3);
or (carry, o1, o2);
endmodule

module multiplier (a, b, m);
input	[31 :0] a;
input	[31 :0] b;
output	[63 :0] m;

wire	[1023 :1]	pp;
wire	[30 :0]	r1c;
wire	[30 :1]	r1s;
wire	[30 :0]	r2c;
wire	[30 :1]	r2s;
wire	[30 :0]	r3c;
wire	[30 :1]	r3s;
wire	[30 :0]	r4c;
wire	[30 :1]	r4s;
wire	[30 :0]	r5c;
wire	[30 :1]	r5s;
wire	[30 :0]	r6c;
wire	[30 :1]	r6s;
wire	[30 :0]	r7c;
wire	[30 :1]	r7s;
wire	[30 :0]	r8c;
wire	[30 :1]	r8s;
wire	[30 :0]	r9c;
wire	[30 :1]	r9s;
wire	[30 :0]	r10c;
wire	[30 :1]	r10s;
wire	[30 :0]	r11c;
wire	[30 :1]	r11s;
wire	[30 :0]	r12c;
wire	[30 :1]	r12s;
wire	[30 :0]	r13c;
wire	[30 :1]	r13s;
wire	[30 :0]	r14c;
wire	[30 :1]	r14s;
wire	[30 :0]	r15c;
wire	[30 :1]	r15s;
wire	[30 :0]	r16c;
wire	[30 :1]	r16s;
wire	[30 :0]	r17c;
wire	[30 :1]	r17s;
wire	[30 :0]	r18c;
wire	[30 :1]	r18s;
wire	[30 :0]	r19c;
wire	[30 :1]	r19s;
wire	[30 :0]	r20c;
wire	[30 :1]	r20s;
wire	[30 :0]	r21c;
wire	[30 :1]	r21s;
wire	[30 :0]	r22c;
wire	[30 :1]	r22s;
wire	[30 :0]	r23c;
wire	[30 :1]	r23s;
wire	[30 :0]	r24c;
wire	[30 :1]	r24s;
wire	[30 :0]	r25c;
wire	[30 :1]	r25s;
wire	[30 :0]	r26c;
wire	[30 :1]	r26s;
wire	[30 :0]	r27c;
wire	[30 :1]	r27s;
wire	[30 :0]	r28c;
wire	[30 :1]	r28s;
wire	[30 :0]	r29c;
wire	[30 :1]	r29s;
wire	[30 :0]	r30c;
wire	[30 :1]	r30s;
wire	[30 :0]	r31c;
wire	[30 :1]	r31s;
wire	[29 :0]	r32c;

and	(m[0], a[0], b[0]);
and	(pp[1], a[0], b[1]);
and	(pp[2], a[0], b[2]);
and	(pp[3], a[0], b[3]);
and	(pp[4], a[0], b[4]);
and	(pp[5], a[0], b[5]);
and	(pp[6], a[0], b[6]);
and	(pp[7], a[0], b[7]);
and	(pp[8], a[0], b[8]);
and	(pp[9], a[0], b[9]);
and	(pp[10], a[0], b[10]);
and	(pp[11], a[0], b[11]);
and	(pp[12], a[0], b[12]);
and	(pp[13], a[0], b[13]);
and	(pp[14], a[0], b[14]);
and	(pp[15], a[0], b[15]);
and	(pp[16], a[0], b[16]);
and	(pp[17], a[0], b[17]);
and	(pp[18], a[0], b[18]);
and	(pp[19], a[0], b[19]);
and	(pp[20], a[0], b[20]);
and	(pp[21], a[0], b[21]);
and	(pp[22], a[0], b[22]);
and	(pp[23], a[0], b[23]);
and	(pp[24], a[0], b[24]);
and	(pp[25], a[0], b[25]);
and	(pp[26], a[0], b[26]);
and	(pp[27], a[0], b[27]);
and	(pp[28], a[0], b[28]);
and	(pp[29], a[0], b[29]);
and	(pp[30], a[0], b[30]);
and	(pp[31], a[0], b[31]);
and	(pp[32], a[1], b[0]);
and	(pp[33], a[1], b[1]);
and	(pp[34], a[1], b[2]);
and	(pp[35], a[1], b[3]);
and	(pp[36], a[1], b[4]);
and	(pp[37], a[1], b[5]);
and	(pp[38], a[1], b[6]);
and	(pp[39], a[1], b[7]);
and	(pp[40], a[1], b[8]);
and	(pp[41], a[1], b[9]);
and	(pp[42], a[1], b[10]);
and	(pp[43], a[1], b[11]);
and	(pp[44], a[1], b[12]);
and	(pp[45], a[1], b[13]);
and	(pp[46], a[1], b[14]);
and	(pp[47], a[1], b[15]);
and	(pp[48], a[1], b[16]);
and	(pp[49], a[1], b[17]);
and	(pp[50], a[1], b[18]);
and	(pp[51], a[1], b[19]);
and	(pp[52], a[1], b[20]);
and	(pp[53], a[1], b[21]);
and	(pp[54], a[1], b[22]);
and	(pp[55], a[1], b[23]);
and	(pp[56], a[1], b[24]);
and	(pp[57], a[1], b[25]);
and	(pp[58], a[1], b[26]);
and	(pp[59], a[1], b[27]);
and	(pp[60], a[1], b[28]);
and	(pp[61], a[1], b[29]);
and	(pp[62], a[1], b[30]);
and	(pp[63], a[1], b[31]);
and	(pp[64], a[2], b[0]);
and	(pp[65], a[2], b[1]);
and	(pp[66], a[2], b[2]);
and	(pp[67], a[2], b[3]);
and	(pp[68], a[2], b[4]);
and	(pp[69], a[2], b[5]);
and	(pp[70], a[2], b[6]);
and	(pp[71], a[2], b[7]);
and	(pp[72], a[2], b[8]);
and	(pp[73], a[2], b[9]);
and	(pp[74], a[2], b[10]);
and	(pp[75], a[2], b[11]);
and	(pp[76], a[2], b[12]);
and	(pp[77], a[2], b[13]);
and	(pp[78], a[2], b[14]);
and	(pp[79], a[2], b[15]);
and	(pp[80], a[2], b[16]);
and	(pp[81], a[2], b[17]);
and	(pp[82], a[2], b[18]);
and	(pp[83], a[2], b[19]);
and	(pp[84], a[2], b[20]);
and	(pp[85], a[2], b[21]);
and	(pp[86], a[2], b[22]);
and	(pp[87], a[2], b[23]);
and	(pp[88], a[2], b[24]);
and	(pp[89], a[2], b[25]);
and	(pp[90], a[2], b[26]);
and	(pp[91], a[2], b[27]);
and	(pp[92], a[2], b[28]);
and	(pp[93], a[2], b[29]);
and	(pp[94], a[2], b[30]);
and	(pp[95], a[2], b[31]);
and	(pp[96], a[3], b[0]);
and	(pp[97], a[3], b[1]);
and	(pp[98], a[3], b[2]);
and	(pp[99], a[3], b[3]);
and	(pp[100], a[3], b[4]);
and	(pp[101], a[3], b[5]);
and	(pp[102], a[3], b[6]);
and	(pp[103], a[3], b[7]);
and	(pp[104], a[3], b[8]);
and	(pp[105], a[3], b[9]);
and	(pp[106], a[3], b[10]);
and	(pp[107], a[3], b[11]);
and	(pp[108], a[3], b[12]);
and	(pp[109], a[3], b[13]);
and	(pp[110], a[3], b[14]);
and	(pp[111], a[3], b[15]);
and	(pp[112], a[3], b[16]);
and	(pp[113], a[3], b[17]);
and	(pp[114], a[3], b[18]);
and	(pp[115], a[3], b[19]);
and	(pp[116], a[3], b[20]);
and	(pp[117], a[3], b[21]);
and	(pp[118], a[3], b[22]);
and	(pp[119], a[3], b[23]);
and	(pp[120], a[3], b[24]);
and	(pp[121], a[3], b[25]);
and	(pp[122], a[3], b[26]);
and	(pp[123], a[3], b[27]);
and	(pp[124], a[3], b[28]);
and	(pp[125], a[3], b[29]);
and	(pp[126], a[3], b[30]);
and	(pp[127], a[3], b[31]);
and	(pp[128], a[4], b[0]);
and	(pp[129], a[4], b[1]);
and	(pp[130], a[4], b[2]);
and	(pp[131], a[4], b[3]);
and	(pp[132], a[4], b[4]);
and	(pp[133], a[4], b[5]);
and	(pp[134], a[4], b[6]);
and	(pp[135], a[4], b[7]);
and	(pp[136], a[4], b[8]);
and	(pp[137], a[4], b[9]);
and	(pp[138], a[4], b[10]);
and	(pp[139], a[4], b[11]);
and	(pp[140], a[4], b[12]);
and	(pp[141], a[4], b[13]);
and	(pp[142], a[4], b[14]);
and	(pp[143], a[4], b[15]);
and	(pp[144], a[4], b[16]);
and	(pp[145], a[4], b[17]);
and	(pp[146], a[4], b[18]);
and	(pp[147], a[4], b[19]);
and	(pp[148], a[4], b[20]);
and	(pp[149], a[4], b[21]);
and	(pp[150], a[4], b[22]);
and	(pp[151], a[4], b[23]);
and	(pp[152], a[4], b[24]);
and	(pp[153], a[4], b[25]);
and	(pp[154], a[4], b[26]);
and	(pp[155], a[4], b[27]);
and	(pp[156], a[4], b[28]);
and	(pp[157], a[4], b[29]);
and	(pp[158], a[4], b[30]);
and	(pp[159], a[4], b[31]);
and	(pp[160], a[5], b[0]);
and	(pp[161], a[5], b[1]);
and	(pp[162], a[5], b[2]);
and	(pp[163], a[5], b[3]);
and	(pp[164], a[5], b[4]);
and	(pp[165], a[5], b[5]);
and	(pp[166], a[5], b[6]);
and	(pp[167], a[5], b[7]);
and	(pp[168], a[5], b[8]);
and	(pp[169], a[5], b[9]);
and	(pp[170], a[5], b[10]);
and	(pp[171], a[5], b[11]);
and	(pp[172], a[5], b[12]);
and	(pp[173], a[5], b[13]);
and	(pp[174], a[5], b[14]);
and	(pp[175], a[5], b[15]);
and	(pp[176], a[5], b[16]);
and	(pp[177], a[5], b[17]);
and	(pp[178], a[5], b[18]);
and	(pp[179], a[5], b[19]);
and	(pp[180], a[5], b[20]);
and	(pp[181], a[5], b[21]);
and	(pp[182], a[5], b[22]);
and	(pp[183], a[5], b[23]);
and	(pp[184], a[5], b[24]);
and	(pp[185], a[5], b[25]);
and	(pp[186], a[5], b[26]);
and	(pp[187], a[5], b[27]);
and	(pp[188], a[5], b[28]);
and	(pp[189], a[5], b[29]);
and	(pp[190], a[5], b[30]);
and	(pp[191], a[5], b[31]);
and	(pp[192], a[6], b[0]);
and	(pp[193], a[6], b[1]);
and	(pp[194], a[6], b[2]);
and	(pp[195], a[6], b[3]);
and	(pp[196], a[6], b[4]);
and	(pp[197], a[6], b[5]);
and	(pp[198], a[6], b[6]);
and	(pp[199], a[6], b[7]);
and	(pp[200], a[6], b[8]);
and	(pp[201], a[6], b[9]);
and	(pp[202], a[6], b[10]);
and	(pp[203], a[6], b[11]);
and	(pp[204], a[6], b[12]);
and	(pp[205], a[6], b[13]);
and	(pp[206], a[6], b[14]);
and	(pp[207], a[6], b[15]);
and	(pp[208], a[6], b[16]);
and	(pp[209], a[6], b[17]);
and	(pp[210], a[6], b[18]);
and	(pp[211], a[6], b[19]);
and	(pp[212], a[6], b[20]);
and	(pp[213], a[6], b[21]);
and	(pp[214], a[6], b[22]);
and	(pp[215], a[6], b[23]);
and	(pp[216], a[6], b[24]);
and	(pp[217], a[6], b[25]);
and	(pp[218], a[6], b[26]);
and	(pp[219], a[6], b[27]);
and	(pp[220], a[6], b[28]);
and	(pp[221], a[6], b[29]);
and	(pp[222], a[6], b[30]);
and	(pp[223], a[6], b[31]);
and	(pp[224], a[7], b[0]);
and	(pp[225], a[7], b[1]);
and	(pp[226], a[7], b[2]);
and	(pp[227], a[7], b[3]);
and	(pp[228], a[7], b[4]);
and	(pp[229], a[7], b[5]);
and	(pp[230], a[7], b[6]);
and	(pp[231], a[7], b[7]);
and	(pp[232], a[7], b[8]);
and	(pp[233], a[7], b[9]);
and	(pp[234], a[7], b[10]);
and	(pp[235], a[7], b[11]);
and	(pp[236], a[7], b[12]);
and	(pp[237], a[7], b[13]);
and	(pp[238], a[7], b[14]);
and	(pp[239], a[7], b[15]);
and	(pp[240], a[7], b[16]);
and	(pp[241], a[7], b[17]);
and	(pp[242], a[7], b[18]);
and	(pp[243], a[7], b[19]);
and	(pp[244], a[7], b[20]);
and	(pp[245], a[7], b[21]);
and	(pp[246], a[7], b[22]);
and	(pp[247], a[7], b[23]);
and	(pp[248], a[7], b[24]);
and	(pp[249], a[7], b[25]);
and	(pp[250], a[7], b[26]);
and	(pp[251], a[7], b[27]);
and	(pp[252], a[7], b[28]);
and	(pp[253], a[7], b[29]);
and	(pp[254], a[7], b[30]);
and	(pp[255], a[7], b[31]);
and	(pp[256], a[8], b[0]);
and	(pp[257], a[8], b[1]);
and	(pp[258], a[8], b[2]);
and	(pp[259], a[8], b[3]);
and	(pp[260], a[8], b[4]);
and	(pp[261], a[8], b[5]);
and	(pp[262], a[8], b[6]);
and	(pp[263], a[8], b[7]);
and	(pp[264], a[8], b[8]);
and	(pp[265], a[8], b[9]);
and	(pp[266], a[8], b[10]);
and	(pp[267], a[8], b[11]);
and	(pp[268], a[8], b[12]);
and	(pp[269], a[8], b[13]);
and	(pp[270], a[8], b[14]);
and	(pp[271], a[8], b[15]);
and	(pp[272], a[8], b[16]);
and	(pp[273], a[8], b[17]);
and	(pp[274], a[8], b[18]);
and	(pp[275], a[8], b[19]);
and	(pp[276], a[8], b[20]);
and	(pp[277], a[8], b[21]);
and	(pp[278], a[8], b[22]);
and	(pp[279], a[8], b[23]);
and	(pp[280], a[8], b[24]);
and	(pp[281], a[8], b[25]);
and	(pp[282], a[8], b[26]);
and	(pp[283], a[8], b[27]);
and	(pp[284], a[8], b[28]);
and	(pp[285], a[8], b[29]);
and	(pp[286], a[8], b[30]);
and	(pp[287], a[8], b[31]);
and	(pp[288], a[9], b[0]);
and	(pp[289], a[9], b[1]);
and	(pp[290], a[9], b[2]);
and	(pp[291], a[9], b[3]);
and	(pp[292], a[9], b[4]);
and	(pp[293], a[9], b[5]);
and	(pp[294], a[9], b[6]);
and	(pp[295], a[9], b[7]);
and	(pp[296], a[9], b[8]);
and	(pp[297], a[9], b[9]);
and	(pp[298], a[9], b[10]);
and	(pp[299], a[9], b[11]);
and	(pp[300], a[9], b[12]);
and	(pp[301], a[9], b[13]);
and	(pp[302], a[9], b[14]);
and	(pp[303], a[9], b[15]);
and	(pp[304], a[9], b[16]);
and	(pp[305], a[9], b[17]);
and	(pp[306], a[9], b[18]);
and	(pp[307], a[9], b[19]);
and	(pp[308], a[9], b[20]);
and	(pp[309], a[9], b[21]);
and	(pp[310], a[9], b[22]);
and	(pp[311], a[9], b[23]);
and	(pp[312], a[9], b[24]);
and	(pp[313], a[9], b[25]);
and	(pp[314], a[9], b[26]);
and	(pp[315], a[9], b[27]);
and	(pp[316], a[9], b[28]);
and	(pp[317], a[9], b[29]);
and	(pp[318], a[9], b[30]);
and	(pp[319], a[9], b[31]);
and	(pp[320], a[10], b[0]);
and	(pp[321], a[10], b[1]);
and	(pp[322], a[10], b[2]);
and	(pp[323], a[10], b[3]);
and	(pp[324], a[10], b[4]);
and	(pp[325], a[10], b[5]);
and	(pp[326], a[10], b[6]);
and	(pp[327], a[10], b[7]);
and	(pp[328], a[10], b[8]);
and	(pp[329], a[10], b[9]);
and	(pp[330], a[10], b[10]);
and	(pp[331], a[10], b[11]);
and	(pp[332], a[10], b[12]);
and	(pp[333], a[10], b[13]);
and	(pp[334], a[10], b[14]);
and	(pp[335], a[10], b[15]);
and	(pp[336], a[10], b[16]);
and	(pp[337], a[10], b[17]);
and	(pp[338], a[10], b[18]);
and	(pp[339], a[10], b[19]);
and	(pp[340], a[10], b[20]);
and	(pp[341], a[10], b[21]);
and	(pp[342], a[10], b[22]);
and	(pp[343], a[10], b[23]);
and	(pp[344], a[10], b[24]);
and	(pp[345], a[10], b[25]);
and	(pp[346], a[10], b[26]);
and	(pp[347], a[10], b[27]);
and	(pp[348], a[10], b[28]);
and	(pp[349], a[10], b[29]);
and	(pp[350], a[10], b[30]);
and	(pp[351], a[10], b[31]);
and	(pp[352], a[11], b[0]);
and	(pp[353], a[11], b[1]);
and	(pp[354], a[11], b[2]);
and	(pp[355], a[11], b[3]);
and	(pp[356], a[11], b[4]);
and	(pp[357], a[11], b[5]);
and	(pp[358], a[11], b[6]);
and	(pp[359], a[11], b[7]);
and	(pp[360], a[11], b[8]);
and	(pp[361], a[11], b[9]);
and	(pp[362], a[11], b[10]);
and	(pp[363], a[11], b[11]);
and	(pp[364], a[11], b[12]);
and	(pp[365], a[11], b[13]);
and	(pp[366], a[11], b[14]);
and	(pp[367], a[11], b[15]);
and	(pp[368], a[11], b[16]);
and	(pp[369], a[11], b[17]);
and	(pp[370], a[11], b[18]);
and	(pp[371], a[11], b[19]);
and	(pp[372], a[11], b[20]);
and	(pp[373], a[11], b[21]);
and	(pp[374], a[11], b[22]);
and	(pp[375], a[11], b[23]);
and	(pp[376], a[11], b[24]);
and	(pp[377], a[11], b[25]);
and	(pp[378], a[11], b[26]);
and	(pp[379], a[11], b[27]);
and	(pp[380], a[11], b[28]);
and	(pp[381], a[11], b[29]);
and	(pp[382], a[11], b[30]);
and	(pp[383], a[11], b[31]);
and	(pp[384], a[12], b[0]);
and	(pp[385], a[12], b[1]);
and	(pp[386], a[12], b[2]);
and	(pp[387], a[12], b[3]);
and	(pp[388], a[12], b[4]);
and	(pp[389], a[12], b[5]);
and	(pp[390], a[12], b[6]);
and	(pp[391], a[12], b[7]);
and	(pp[392], a[12], b[8]);
and	(pp[393], a[12], b[9]);
and	(pp[394], a[12], b[10]);
and	(pp[395], a[12], b[11]);
and	(pp[396], a[12], b[12]);
and	(pp[397], a[12], b[13]);
and	(pp[398], a[12], b[14]);
and	(pp[399], a[12], b[15]);
and	(pp[400], a[12], b[16]);
and	(pp[401], a[12], b[17]);
and	(pp[402], a[12], b[18]);
and	(pp[403], a[12], b[19]);
and	(pp[404], a[12], b[20]);
and	(pp[405], a[12], b[21]);
and	(pp[406], a[12], b[22]);
and	(pp[407], a[12], b[23]);
and	(pp[408], a[12], b[24]);
and	(pp[409], a[12], b[25]);
and	(pp[410], a[12], b[26]);
and	(pp[411], a[12], b[27]);
and	(pp[412], a[12], b[28]);
and	(pp[413], a[12], b[29]);
and	(pp[414], a[12], b[30]);
and	(pp[415], a[12], b[31]);
and	(pp[416], a[13], b[0]);
and	(pp[417], a[13], b[1]);
and	(pp[418], a[13], b[2]);
and	(pp[419], a[13], b[3]);
and	(pp[420], a[13], b[4]);
and	(pp[421], a[13], b[5]);
and	(pp[422], a[13], b[6]);
and	(pp[423], a[13], b[7]);
and	(pp[424], a[13], b[8]);
and	(pp[425], a[13], b[9]);
and	(pp[426], a[13], b[10]);
and	(pp[427], a[13], b[11]);
and	(pp[428], a[13], b[12]);
and	(pp[429], a[13], b[13]);
and	(pp[430], a[13], b[14]);
and	(pp[431], a[13], b[15]);
and	(pp[432], a[13], b[16]);
and	(pp[433], a[13], b[17]);
and	(pp[434], a[13], b[18]);
and	(pp[435], a[13], b[19]);
and	(pp[436], a[13], b[20]);
and	(pp[437], a[13], b[21]);
and	(pp[438], a[13], b[22]);
and	(pp[439], a[13], b[23]);
and	(pp[440], a[13], b[24]);
and	(pp[441], a[13], b[25]);
and	(pp[442], a[13], b[26]);
and	(pp[443], a[13], b[27]);
and	(pp[444], a[13], b[28]);
and	(pp[445], a[13], b[29]);
and	(pp[446], a[13], b[30]);
and	(pp[447], a[13], b[31]);
and	(pp[448], a[14], b[0]);
and	(pp[449], a[14], b[1]);
and	(pp[450], a[14], b[2]);
and	(pp[451], a[14], b[3]);
and	(pp[452], a[14], b[4]);
and	(pp[453], a[14], b[5]);
and	(pp[454], a[14], b[6]);
and	(pp[455], a[14], b[7]);
and	(pp[456], a[14], b[8]);
and	(pp[457], a[14], b[9]);
and	(pp[458], a[14], b[10]);
and	(pp[459], a[14], b[11]);
and	(pp[460], a[14], b[12]);
and	(pp[461], a[14], b[13]);
and	(pp[462], a[14], b[14]);
and	(pp[463], a[14], b[15]);
and	(pp[464], a[14], b[16]);
and	(pp[465], a[14], b[17]);
and	(pp[466], a[14], b[18]);
and	(pp[467], a[14], b[19]);
and	(pp[468], a[14], b[20]);
and	(pp[469], a[14], b[21]);
and	(pp[470], a[14], b[22]);
and	(pp[471], a[14], b[23]);
and	(pp[472], a[14], b[24]);
and	(pp[473], a[14], b[25]);
and	(pp[474], a[14], b[26]);
and	(pp[475], a[14], b[27]);
and	(pp[476], a[14], b[28]);
and	(pp[477], a[14], b[29]);
and	(pp[478], a[14], b[30]);
and	(pp[479], a[14], b[31]);
and	(pp[480], a[15], b[0]);
and	(pp[481], a[15], b[1]);
and	(pp[482], a[15], b[2]);
and	(pp[483], a[15], b[3]);
and	(pp[484], a[15], b[4]);
and	(pp[485], a[15], b[5]);
and	(pp[486], a[15], b[6]);
and	(pp[487], a[15], b[7]);
and	(pp[488], a[15], b[8]);
and	(pp[489], a[15], b[9]);
and	(pp[490], a[15], b[10]);
and	(pp[491], a[15], b[11]);
and	(pp[492], a[15], b[12]);
and	(pp[493], a[15], b[13]);
and	(pp[494], a[15], b[14]);
and	(pp[495], a[15], b[15]);
and	(pp[496], a[15], b[16]);
and	(pp[497], a[15], b[17]);
and	(pp[498], a[15], b[18]);
and	(pp[499], a[15], b[19]);
and	(pp[500], a[15], b[20]);
and	(pp[501], a[15], b[21]);
and	(pp[502], a[15], b[22]);
and	(pp[503], a[15], b[23]);
and	(pp[504], a[15], b[24]);
and	(pp[505], a[15], b[25]);
and	(pp[506], a[15], b[26]);
and	(pp[507], a[15], b[27]);
and	(pp[508], a[15], b[28]);
and	(pp[509], a[15], b[29]);
and	(pp[510], a[15], b[30]);
and	(pp[511], a[15], b[31]);
and	(pp[512], a[16], b[0]);
and	(pp[513], a[16], b[1]);
and	(pp[514], a[16], b[2]);
and	(pp[515], a[16], b[3]);
and	(pp[516], a[16], b[4]);
and	(pp[517], a[16], b[5]);
and	(pp[518], a[16], b[6]);
and	(pp[519], a[16], b[7]);
and	(pp[520], a[16], b[8]);
and	(pp[521], a[16], b[9]);
and	(pp[522], a[16], b[10]);
and	(pp[523], a[16], b[11]);
and	(pp[524], a[16], b[12]);
and	(pp[525], a[16], b[13]);
and	(pp[526], a[16], b[14]);
and	(pp[527], a[16], b[15]);
and	(pp[528], a[16], b[16]);
and	(pp[529], a[16], b[17]);
and	(pp[530], a[16], b[18]);
and	(pp[531], a[16], b[19]);
and	(pp[532], a[16], b[20]);
and	(pp[533], a[16], b[21]);
and	(pp[534], a[16], b[22]);
and	(pp[535], a[16], b[23]);
and	(pp[536], a[16], b[24]);
and	(pp[537], a[16], b[25]);
and	(pp[538], a[16], b[26]);
and	(pp[539], a[16], b[27]);
and	(pp[540], a[16], b[28]);
and	(pp[541], a[16], b[29]);
and	(pp[542], a[16], b[30]);
and	(pp[543], a[16], b[31]);
and	(pp[544], a[17], b[0]);
and	(pp[545], a[17], b[1]);
and	(pp[546], a[17], b[2]);
and	(pp[547], a[17], b[3]);
and	(pp[548], a[17], b[4]);
and	(pp[549], a[17], b[5]);
and	(pp[550], a[17], b[6]);
and	(pp[551], a[17], b[7]);
and	(pp[552], a[17], b[8]);
and	(pp[553], a[17], b[9]);
and	(pp[554], a[17], b[10]);
and	(pp[555], a[17], b[11]);
and	(pp[556], a[17], b[12]);
and	(pp[557], a[17], b[13]);
and	(pp[558], a[17], b[14]);
and	(pp[559], a[17], b[15]);
and	(pp[560], a[17], b[16]);
and	(pp[561], a[17], b[17]);
and	(pp[562], a[17], b[18]);
and	(pp[563], a[17], b[19]);
and	(pp[564], a[17], b[20]);
and	(pp[565], a[17], b[21]);
and	(pp[566], a[17], b[22]);
and	(pp[567], a[17], b[23]);
and	(pp[568], a[17], b[24]);
and	(pp[569], a[17], b[25]);
and	(pp[570], a[17], b[26]);
and	(pp[571], a[17], b[27]);
and	(pp[572], a[17], b[28]);
and	(pp[573], a[17], b[29]);
and	(pp[574], a[17], b[30]);
and	(pp[575], a[17], b[31]);
and	(pp[576], a[18], b[0]);
and	(pp[577], a[18], b[1]);
and	(pp[578], a[18], b[2]);
and	(pp[579], a[18], b[3]);
and	(pp[580], a[18], b[4]);
and	(pp[581], a[18], b[5]);
and	(pp[582], a[18], b[6]);
and	(pp[583], a[18], b[7]);
and	(pp[584], a[18], b[8]);
and	(pp[585], a[18], b[9]);
and	(pp[586], a[18], b[10]);
and	(pp[587], a[18], b[11]);
and	(pp[588], a[18], b[12]);
and	(pp[589], a[18], b[13]);
and	(pp[590], a[18], b[14]);
and	(pp[591], a[18], b[15]);
and	(pp[592], a[18], b[16]);
and	(pp[593], a[18], b[17]);
and	(pp[594], a[18], b[18]);
and	(pp[595], a[18], b[19]);
and	(pp[596], a[18], b[20]);
and	(pp[597], a[18], b[21]);
and	(pp[598], a[18], b[22]);
and	(pp[599], a[18], b[23]);
and	(pp[600], a[18], b[24]);
and	(pp[601], a[18], b[25]);
and	(pp[602], a[18], b[26]);
and	(pp[603], a[18], b[27]);
and	(pp[604], a[18], b[28]);
and	(pp[605], a[18], b[29]);
and	(pp[606], a[18], b[30]);
and	(pp[607], a[18], b[31]);
and	(pp[608], a[19], b[0]);
and	(pp[609], a[19], b[1]);
and	(pp[610], a[19], b[2]);
and	(pp[611], a[19], b[3]);
and	(pp[612], a[19], b[4]);
and	(pp[613], a[19], b[5]);
and	(pp[614], a[19], b[6]);
and	(pp[615], a[19], b[7]);
and	(pp[616], a[19], b[8]);
and	(pp[617], a[19], b[9]);
and	(pp[618], a[19], b[10]);
and	(pp[619], a[19], b[11]);
and	(pp[620], a[19], b[12]);
and	(pp[621], a[19], b[13]);
and	(pp[622], a[19], b[14]);
and	(pp[623], a[19], b[15]);
and	(pp[624], a[19], b[16]);
and	(pp[625], a[19], b[17]);
and	(pp[626], a[19], b[18]);
and	(pp[627], a[19], b[19]);
and	(pp[628], a[19], b[20]);
and	(pp[629], a[19], b[21]);
and	(pp[630], a[19], b[22]);
and	(pp[631], a[19], b[23]);
and	(pp[632], a[19], b[24]);
and	(pp[633], a[19], b[25]);
and	(pp[634], a[19], b[26]);
and	(pp[635], a[19], b[27]);
and	(pp[636], a[19], b[28]);
and	(pp[637], a[19], b[29]);
and	(pp[638], a[19], b[30]);
and	(pp[639], a[19], b[31]);
and	(pp[640], a[20], b[0]);
and	(pp[641], a[20], b[1]);
and	(pp[642], a[20], b[2]);
and	(pp[643], a[20], b[3]);
and	(pp[644], a[20], b[4]);
and	(pp[645], a[20], b[5]);
and	(pp[646], a[20], b[6]);
and	(pp[647], a[20], b[7]);
and	(pp[648], a[20], b[8]);
and	(pp[649], a[20], b[9]);
and	(pp[650], a[20], b[10]);
and	(pp[651], a[20], b[11]);
and	(pp[652], a[20], b[12]);
and	(pp[653], a[20], b[13]);
and	(pp[654], a[20], b[14]);
and	(pp[655], a[20], b[15]);
and	(pp[656], a[20], b[16]);
and	(pp[657], a[20], b[17]);
and	(pp[658], a[20], b[18]);
and	(pp[659], a[20], b[19]);
and	(pp[660], a[20], b[20]);
and	(pp[661], a[20], b[21]);
and	(pp[662], a[20], b[22]);
and	(pp[663], a[20], b[23]);
and	(pp[664], a[20], b[24]);
and	(pp[665], a[20], b[25]);
and	(pp[666], a[20], b[26]);
and	(pp[667], a[20], b[27]);
and	(pp[668], a[20], b[28]);
and	(pp[669], a[20], b[29]);
and	(pp[670], a[20], b[30]);
and	(pp[671], a[20], b[31]);
and	(pp[672], a[21], b[0]);
and	(pp[673], a[21], b[1]);
and	(pp[674], a[21], b[2]);
and	(pp[675], a[21], b[3]);
and	(pp[676], a[21], b[4]);
and	(pp[677], a[21], b[5]);
and	(pp[678], a[21], b[6]);
and	(pp[679], a[21], b[7]);
and	(pp[680], a[21], b[8]);
and	(pp[681], a[21], b[9]);
and	(pp[682], a[21], b[10]);
and	(pp[683], a[21], b[11]);
and	(pp[684], a[21], b[12]);
and	(pp[685], a[21], b[13]);
and	(pp[686], a[21], b[14]);
and	(pp[687], a[21], b[15]);
and	(pp[688], a[21], b[16]);
and	(pp[689], a[21], b[17]);
and	(pp[690], a[21], b[18]);
and	(pp[691], a[21], b[19]);
and	(pp[692], a[21], b[20]);
and	(pp[693], a[21], b[21]);
and	(pp[694], a[21], b[22]);
and	(pp[695], a[21], b[23]);
and	(pp[696], a[21], b[24]);
and	(pp[697], a[21], b[25]);
and	(pp[698], a[21], b[26]);
and	(pp[699], a[21], b[27]);
and	(pp[700], a[21], b[28]);
and	(pp[701], a[21], b[29]);
and	(pp[702], a[21], b[30]);
and	(pp[703], a[21], b[31]);
and	(pp[704], a[22], b[0]);
and	(pp[705], a[22], b[1]);
and	(pp[706], a[22], b[2]);
and	(pp[707], a[22], b[3]);
and	(pp[708], a[22], b[4]);
and	(pp[709], a[22], b[5]);
and	(pp[710], a[22], b[6]);
and	(pp[711], a[22], b[7]);
and	(pp[712], a[22], b[8]);
and	(pp[713], a[22], b[9]);
and	(pp[714], a[22], b[10]);
and	(pp[715], a[22], b[11]);
and	(pp[716], a[22], b[12]);
and	(pp[717], a[22], b[13]);
and	(pp[718], a[22], b[14]);
and	(pp[719], a[22], b[15]);
and	(pp[720], a[22], b[16]);
and	(pp[721], a[22], b[17]);
and	(pp[722], a[22], b[18]);
and	(pp[723], a[22], b[19]);
and	(pp[724], a[22], b[20]);
and	(pp[725], a[22], b[21]);
and	(pp[726], a[22], b[22]);
and	(pp[727], a[22], b[23]);
and	(pp[728], a[22], b[24]);
and	(pp[729], a[22], b[25]);
and	(pp[730], a[22], b[26]);
and	(pp[731], a[22], b[27]);
and	(pp[732], a[22], b[28]);
and	(pp[733], a[22], b[29]);
and	(pp[734], a[22], b[30]);
and	(pp[735], a[22], b[31]);
and	(pp[736], a[23], b[0]);
and	(pp[737], a[23], b[1]);
and	(pp[738], a[23], b[2]);
and	(pp[739], a[23], b[3]);
and	(pp[740], a[23], b[4]);
and	(pp[741], a[23], b[5]);
and	(pp[742], a[23], b[6]);
and	(pp[743], a[23], b[7]);
and	(pp[744], a[23], b[8]);
and	(pp[745], a[23], b[9]);
and	(pp[746], a[23], b[10]);
and	(pp[747], a[23], b[11]);
and	(pp[748], a[23], b[12]);
and	(pp[749], a[23], b[13]);
and	(pp[750], a[23], b[14]);
and	(pp[751], a[23], b[15]);
and	(pp[752], a[23], b[16]);
and	(pp[753], a[23], b[17]);
and	(pp[754], a[23], b[18]);
and	(pp[755], a[23], b[19]);
and	(pp[756], a[23], b[20]);
and	(pp[757], a[23], b[21]);
and	(pp[758], a[23], b[22]);
and	(pp[759], a[23], b[23]);
and	(pp[760], a[23], b[24]);
and	(pp[761], a[23], b[25]);
and	(pp[762], a[23], b[26]);
and	(pp[763], a[23], b[27]);
and	(pp[764], a[23], b[28]);
and	(pp[765], a[23], b[29]);
and	(pp[766], a[23], b[30]);
and	(pp[767], a[23], b[31]);
and	(pp[768], a[24], b[0]);
and	(pp[769], a[24], b[1]);
and	(pp[770], a[24], b[2]);
and	(pp[771], a[24], b[3]);
and	(pp[772], a[24], b[4]);
and	(pp[773], a[24], b[5]);
and	(pp[774], a[24], b[6]);
and	(pp[775], a[24], b[7]);
and	(pp[776], a[24], b[8]);
and	(pp[777], a[24], b[9]);
and	(pp[778], a[24], b[10]);
and	(pp[779], a[24], b[11]);
and	(pp[780], a[24], b[12]);
and	(pp[781], a[24], b[13]);
and	(pp[782], a[24], b[14]);
and	(pp[783], a[24], b[15]);
and	(pp[784], a[24], b[16]);
and	(pp[785], a[24], b[17]);
and	(pp[786], a[24], b[18]);
and	(pp[787], a[24], b[19]);
and	(pp[788], a[24], b[20]);
and	(pp[789], a[24], b[21]);
and	(pp[790], a[24], b[22]);
and	(pp[791], a[24], b[23]);
and	(pp[792], a[24], b[24]);
and	(pp[793], a[24], b[25]);
and	(pp[794], a[24], b[26]);
and	(pp[795], a[24], b[27]);
and	(pp[796], a[24], b[28]);
and	(pp[797], a[24], b[29]);
and	(pp[798], a[24], b[30]);
and	(pp[799], a[24], b[31]);
and	(pp[800], a[25], b[0]);
and	(pp[801], a[25], b[1]);
and	(pp[802], a[25], b[2]);
and	(pp[803], a[25], b[3]);
and	(pp[804], a[25], b[4]);
and	(pp[805], a[25], b[5]);
and	(pp[806], a[25], b[6]);
and	(pp[807], a[25], b[7]);
and	(pp[808], a[25], b[8]);
and	(pp[809], a[25], b[9]);
and	(pp[810], a[25], b[10]);
and	(pp[811], a[25], b[11]);
and	(pp[812], a[25], b[12]);
and	(pp[813], a[25], b[13]);
and	(pp[814], a[25], b[14]);
and	(pp[815], a[25], b[15]);
and	(pp[816], a[25], b[16]);
and	(pp[817], a[25], b[17]);
and	(pp[818], a[25], b[18]);
and	(pp[819], a[25], b[19]);
and	(pp[820], a[25], b[20]);
and	(pp[821], a[25], b[21]);
and	(pp[822], a[25], b[22]);
and	(pp[823], a[25], b[23]);
and	(pp[824], a[25], b[24]);
and	(pp[825], a[25], b[25]);
and	(pp[826], a[25], b[26]);
and	(pp[827], a[25], b[27]);
and	(pp[828], a[25], b[28]);
and	(pp[829], a[25], b[29]);
and	(pp[830], a[25], b[30]);
and	(pp[831], a[25], b[31]);
and	(pp[832], a[26], b[0]);
and	(pp[833], a[26], b[1]);
and	(pp[834], a[26], b[2]);
and	(pp[835], a[26], b[3]);
and	(pp[836], a[26], b[4]);
and	(pp[837], a[26], b[5]);
and	(pp[838], a[26], b[6]);
and	(pp[839], a[26], b[7]);
and	(pp[840], a[26], b[8]);
and	(pp[841], a[26], b[9]);
and	(pp[842], a[26], b[10]);
and	(pp[843], a[26], b[11]);
and	(pp[844], a[26], b[12]);
and	(pp[845], a[26], b[13]);
and	(pp[846], a[26], b[14]);
and	(pp[847], a[26], b[15]);
and	(pp[848], a[26], b[16]);
and	(pp[849], a[26], b[17]);
and	(pp[850], a[26], b[18]);
and	(pp[851], a[26], b[19]);
and	(pp[852], a[26], b[20]);
and	(pp[853], a[26], b[21]);
and	(pp[854], a[26], b[22]);
and	(pp[855], a[26], b[23]);
and	(pp[856], a[26], b[24]);
and	(pp[857], a[26], b[25]);
and	(pp[858], a[26], b[26]);
and	(pp[859], a[26], b[27]);
and	(pp[860], a[26], b[28]);
and	(pp[861], a[26], b[29]);
and	(pp[862], a[26], b[30]);
and	(pp[863], a[26], b[31]);
and	(pp[864], a[27], b[0]);
and	(pp[865], a[27], b[1]);
and	(pp[866], a[27], b[2]);
and	(pp[867], a[27], b[3]);
and	(pp[868], a[27], b[4]);
and	(pp[869], a[27], b[5]);
and	(pp[870], a[27], b[6]);
and	(pp[871], a[27], b[7]);
and	(pp[872], a[27], b[8]);
and	(pp[873], a[27], b[9]);
and	(pp[874], a[27], b[10]);
and	(pp[875], a[27], b[11]);
and	(pp[876], a[27], b[12]);
and	(pp[877], a[27], b[13]);
and	(pp[878], a[27], b[14]);
and	(pp[879], a[27], b[15]);
and	(pp[880], a[27], b[16]);
and	(pp[881], a[27], b[17]);
and	(pp[882], a[27], b[18]);
and	(pp[883], a[27], b[19]);
and	(pp[884], a[27], b[20]);
and	(pp[885], a[27], b[21]);
and	(pp[886], a[27], b[22]);
and	(pp[887], a[27], b[23]);
and	(pp[888], a[27], b[24]);
and	(pp[889], a[27], b[25]);
and	(pp[890], a[27], b[26]);
and	(pp[891], a[27], b[27]);
and	(pp[892], a[27], b[28]);
and	(pp[893], a[27], b[29]);
and	(pp[894], a[27], b[30]);
and	(pp[895], a[27], b[31]);
and	(pp[896], a[28], b[0]);
and	(pp[897], a[28], b[1]);
and	(pp[898], a[28], b[2]);
and	(pp[899], a[28], b[3]);
and	(pp[900], a[28], b[4]);
and	(pp[901], a[28], b[5]);
and	(pp[902], a[28], b[6]);
and	(pp[903], a[28], b[7]);
and	(pp[904], a[28], b[8]);
and	(pp[905], a[28], b[9]);
and	(pp[906], a[28], b[10]);
and	(pp[907], a[28], b[11]);
and	(pp[908], a[28], b[12]);
and	(pp[909], a[28], b[13]);
and	(pp[910], a[28], b[14]);
and	(pp[911], a[28], b[15]);
and	(pp[912], a[28], b[16]);
and	(pp[913], a[28], b[17]);
and	(pp[914], a[28], b[18]);
and	(pp[915], a[28], b[19]);
and	(pp[916], a[28], b[20]);
and	(pp[917], a[28], b[21]);
and	(pp[918], a[28], b[22]);
and	(pp[919], a[28], b[23]);
and	(pp[920], a[28], b[24]);
and	(pp[921], a[28], b[25]);
and	(pp[922], a[28], b[26]);
and	(pp[923], a[28], b[27]);
and	(pp[924], a[28], b[28]);
and	(pp[925], a[28], b[29]);
and	(pp[926], a[28], b[30]);
and	(pp[927], a[28], b[31]);
and	(pp[928], a[29], b[0]);
and	(pp[929], a[29], b[1]);
and	(pp[930], a[29], b[2]);
and	(pp[931], a[29], b[3]);
and	(pp[932], a[29], b[4]);
and	(pp[933], a[29], b[5]);
and	(pp[934], a[29], b[6]);
and	(pp[935], a[29], b[7]);
and	(pp[936], a[29], b[8]);
and	(pp[937], a[29], b[9]);
and	(pp[938], a[29], b[10]);
and	(pp[939], a[29], b[11]);
and	(pp[940], a[29], b[12]);
and	(pp[941], a[29], b[13]);
and	(pp[942], a[29], b[14]);
and	(pp[943], a[29], b[15]);
and	(pp[944], a[29], b[16]);
and	(pp[945], a[29], b[17]);
and	(pp[946], a[29], b[18]);
and	(pp[947], a[29], b[19]);
and	(pp[948], a[29], b[20]);
and	(pp[949], a[29], b[21]);
and	(pp[950], a[29], b[22]);
and	(pp[951], a[29], b[23]);
and	(pp[952], a[29], b[24]);
and	(pp[953], a[29], b[25]);
and	(pp[954], a[29], b[26]);
and	(pp[955], a[29], b[27]);
and	(pp[956], a[29], b[28]);
and	(pp[957], a[29], b[29]);
and	(pp[958], a[29], b[30]);
and	(pp[959], a[29], b[31]);
and	(pp[960], a[30], b[0]);
and	(pp[961], a[30], b[1]);
and	(pp[962], a[30], b[2]);
and	(pp[963], a[30], b[3]);
and	(pp[964], a[30], b[4]);
and	(pp[965], a[30], b[5]);
and	(pp[966], a[30], b[6]);
and	(pp[967], a[30], b[7]);
and	(pp[968], a[30], b[8]);
and	(pp[969], a[30], b[9]);
and	(pp[970], a[30], b[10]);
and	(pp[971], a[30], b[11]);
and	(pp[972], a[30], b[12]);
and	(pp[973], a[30], b[13]);
and	(pp[974], a[30], b[14]);
and	(pp[975], a[30], b[15]);
and	(pp[976], a[30], b[16]);
and	(pp[977], a[30], b[17]);
and	(pp[978], a[30], b[18]);
and	(pp[979], a[30], b[19]);
and	(pp[980], a[30], b[20]);
and	(pp[981], a[30], b[21]);
and	(pp[982], a[30], b[22]);
and	(pp[983], a[30], b[23]);
and	(pp[984], a[30], b[24]);
and	(pp[985], a[30], b[25]);
and	(pp[986], a[30], b[26]);
and	(pp[987], a[30], b[27]);
and	(pp[988], a[30], b[28]);
and	(pp[989], a[30], b[29]);
and	(pp[990], a[30], b[30]);
and	(pp[991], a[30], b[31]);
and	(pp[992], a[31], b[0]);
and	(pp[993], a[31], b[1]);
and	(pp[994], a[31], b[2]);
and	(pp[995], a[31], b[3]);
and	(pp[996], a[31], b[4]);
and	(pp[997], a[31], b[5]);
and	(pp[998], a[31], b[6]);
and	(pp[999], a[31], b[7]);
and	(pp[1000], a[31], b[8]);
and	(pp[1001], a[31], b[9]);
and	(pp[1002], a[31], b[10]);
and	(pp[1003], a[31], b[11]);
and	(pp[1004], a[31], b[12]);
and	(pp[1005], a[31], b[13]);
and	(pp[1006], a[31], b[14]);
and	(pp[1007], a[31], b[15]);
and	(pp[1008], a[31], b[16]);
and	(pp[1009], a[31], b[17]);
and	(pp[1010], a[31], b[18]);
and	(pp[1011], a[31], b[19]);
and	(pp[1012], a[31], b[20]);
and	(pp[1013], a[31], b[21]);
and	(pp[1014], a[31], b[22]);
and	(pp[1015], a[31], b[23]);
and	(pp[1016], a[31], b[24]);
and	(pp[1017], a[31], b[25]);
and	(pp[1018], a[31], b[26]);
and	(pp[1019], a[31], b[27]);
and	(pp[1020], a[31], b[28]);
and	(pp[1021], a[31], b[29]);
and	(pp[1022], a[31], b[30]);
and	(pp[1023], a[31], b[31]);

HA	inst1025	(pp[32], pp[1], m[1], r1c[0]);
FA	inst1026	(pp[33], pp[2], r1c[0], r1s[1], r1c[1]);
FA	inst1027	(pp[34], pp[3], r1c[1], r1s[2], r1c[2]);
FA	inst1028	(pp[35], pp[4], r1c[2], r1s[3], r1c[3]);
FA	inst1029	(pp[36], pp[5], r1c[3], r1s[4], r1c[4]);
FA	inst1030	(pp[37], pp[6], r1c[4], r1s[5], r1c[5]);
FA	inst1031	(pp[38], pp[7], r1c[5], r1s[6], r1c[6]);
FA	inst1032	(pp[39], pp[8], r1c[6], r1s[7], r1c[7]);
FA	inst1033	(pp[40], pp[9], r1c[7], r1s[8], r1c[8]);
FA	inst1034	(pp[41], pp[10], r1c[8], r1s[9], r1c[9]);
FA	inst1035	(pp[42], pp[11], r1c[9], r1s[10], r1c[10]);
FA	inst1036	(pp[43], pp[12], r1c[10], r1s[11], r1c[11]);
FA	inst1037	(pp[44], pp[13], r1c[11], r1s[12], r1c[12]);
FA	inst1038	(pp[45], pp[14], r1c[12], r1s[13], r1c[13]);
FA	inst1039	(pp[46], pp[15], r1c[13], r1s[14], r1c[14]);
FA	inst1040	(pp[47], pp[16], r1c[14], r1s[15], r1c[15]);
FA	inst1041	(pp[48], pp[17], r1c[15], r1s[16], r1c[16]);
FA	inst1042	(pp[49], pp[18], r1c[16], r1s[17], r1c[17]);
FA	inst1043	(pp[50], pp[19], r1c[17], r1s[18], r1c[18]);
FA	inst1044	(pp[51], pp[20], r1c[18], r1s[19], r1c[19]);
FA	inst1045	(pp[52], pp[21], r1c[19], r1s[20], r1c[20]);
FA	inst1046	(pp[53], pp[22], r1c[20], r1s[21], r1c[21]);
FA	inst1047	(pp[54], pp[23], r1c[21], r1s[22], r1c[22]);
FA	inst1048	(pp[55], pp[24], r1c[22], r1s[23], r1c[23]);
FA	inst1049	(pp[56], pp[25], r1c[23], r1s[24], r1c[24]);
FA	inst1050	(pp[57], pp[26], r1c[24], r1s[25], r1c[25]);
FA	inst1051	(pp[58], pp[27], r1c[25], r1s[26], r1c[26]);
FA	inst1052	(pp[59], pp[28], r1c[26], r1s[27], r1c[27]);
FA	inst1053	(pp[60], pp[29], r1c[27], r1s[28], r1c[28]);
FA	inst1054	(pp[61], pp[30], r1c[28], r1s[29], r1c[29]);
FA	inst1055	(pp[62], pp[31], r1c[29], r1s[30], r1c[30]);

HA	inst1056	(r1s[1], pp[64], m[2], r2c[0]);
FA	inst1057	(r1s[2], pp[65], r2c[0], r2s[1], r2c[1]);
FA	inst1058	(r1s[3], pp[66], r2c[1], r2s[2], r2c[2]);
FA	inst1059	(r1s[4], pp[67], r2c[2], r2s[3], r2c[3]);
FA	inst1060	(r1s[5], pp[68], r2c[3], r2s[4], r2c[4]);
FA	inst1061	(r1s[6], pp[69], r2c[4], r2s[5], r2c[5]);
FA	inst1062	(r1s[7], pp[70], r2c[5], r2s[6], r2c[6]);
FA	inst1063	(r1s[8], pp[71], r2c[6], r2s[7], r2c[7]);
FA	inst1064	(r1s[9], pp[72], r2c[7], r2s[8], r2c[8]);
FA	inst1065	(r1s[10], pp[73], r2c[8], r2s[9], r2c[9]);
FA	inst1066	(r1s[11], pp[74], r2c[9], r2s[10], r2c[10]);
FA	inst1067	(r1s[12], pp[75], r2c[10], r2s[11], r2c[11]);
FA	inst1068	(r1s[13], pp[76], r2c[11], r2s[12], r2c[12]);
FA	inst1069	(r1s[14], pp[77], r2c[12], r2s[13], r2c[13]);
FA	inst1070	(r1s[15], pp[78], r2c[13], r2s[14], r2c[14]);
FA	inst1071	(r1s[16], pp[79], r2c[14], r2s[15], r2c[15]);
FA	inst1072	(r1s[17], pp[80], r2c[15], r2s[16], r2c[16]);
FA	inst1073	(r1s[18], pp[81], r2c[16], r2s[17], r2c[17]);
FA	inst1074	(r1s[19], pp[82], r2c[17], r2s[18], r2c[18]);
FA	inst1075	(r1s[20], pp[83], r2c[18], r2s[19], r2c[19]);
FA	inst1076	(r1s[21], pp[84], r2c[19], r2s[20], r2c[20]);
FA	inst1077	(r1s[22], pp[85], r2c[20], r2s[21], r2c[21]);
FA	inst1078	(r1s[23], pp[86], r2c[21], r2s[22], r2c[22]);
FA	inst1079	(r1s[24], pp[87], r2c[22], r2s[23], r2c[23]);
FA	inst1080	(r1s[25], pp[88], r2c[23], r2s[24], r2c[24]);
FA	inst1081	(r1s[26], pp[89], r2c[24], r2s[25], r2c[25]);
FA	inst1082	(r1s[27], pp[90], r2c[25], r2s[26], r2c[26]);
FA	inst1083	(r1s[28], pp[91], r2c[26], r2s[27], r2c[27]);
FA	inst1084	(r1s[29], pp[92], r2c[27], r2s[28], r2c[28]);
FA	inst1085	(r1s[30], pp[93], r2c[28], r2s[29], r2c[29]);
FA	inst1086	(r1c[30], pp[63], r2c[29], r2s[30], r2c[30]);

HA	inst1087	(r2s[1], pp[96], m[3], r3c[0]);
FA	inst1088	(r2s[2], pp[97], r3c[0], r3s[1], r3c[1]);
FA	inst1089	(r2s[3], pp[98], r3c[1], r3s[2], r3c[2]);
FA	inst1090	(r2s[4], pp[99], r3c[2], r3s[3], r3c[3]);
FA	inst1091	(r2s[5], pp[100], r3c[3], r3s[4], r3c[4]);
FA	inst1092	(r2s[6], pp[101], r3c[4], r3s[5], r3c[5]);
FA	inst1093	(r2s[7], pp[102], r3c[5], r3s[6], r3c[6]);
FA	inst1094	(r2s[8], pp[103], r3c[6], r3s[7], r3c[7]);
FA	inst1095	(r2s[9], pp[104], r3c[7], r3s[8], r3c[8]);
FA	inst1096	(r2s[10], pp[105], r3c[8], r3s[9], r3c[9]);
FA	inst1097	(r2s[11], pp[106], r3c[9], r3s[10], r3c[10]);
FA	inst1098	(r2s[12], pp[107], r3c[10], r3s[11], r3c[11]);
FA	inst1099	(r2s[13], pp[108], r3c[11], r3s[12], r3c[12]);
FA	inst1100	(r2s[14], pp[109], r3c[12], r3s[13], r3c[13]);
FA	inst1101	(r2s[15], pp[110], r3c[13], r3s[14], r3c[14]);
FA	inst1102	(r2s[16], pp[111], r3c[14], r3s[15], r3c[15]);
FA	inst1103	(r2s[17], pp[112], r3c[15], r3s[16], r3c[16]);
FA	inst1104	(r2s[18], pp[113], r3c[16], r3s[17], r3c[17]);
FA	inst1105	(r2s[19], pp[114], r3c[17], r3s[18], r3c[18]);
FA	inst1106	(r2s[20], pp[115], r3c[18], r3s[19], r3c[19]);
FA	inst1107	(r2s[21], pp[116], r3c[19], r3s[20], r3c[20]);
FA	inst1108	(r2s[22], pp[117], r3c[20], r3s[21], r3c[21]);
FA	inst1109	(r2s[23], pp[118], r3c[21], r3s[22], r3c[22]);
FA	inst1110	(r2s[24], pp[119], r3c[22], r3s[23], r3c[23]);
FA	inst1111	(r2s[25], pp[120], r3c[23], r3s[24], r3c[24]);
FA	inst1112	(r2s[26], pp[121], r3c[24], r3s[25], r3c[25]);
FA	inst1113	(r2s[27], pp[122], r3c[25], r3s[26], r3c[26]);
FA	inst1114	(r2s[28], pp[123], r3c[26], r3s[27], r3c[27]);
FA	inst1115	(r2s[29], pp[124], r3c[27], r3s[28], r3c[28]);
FA	inst1116	(r2s[30], pp[94], r3c[28], r3s[29], r3c[29]);
FA	inst1117	(r2c[30], pp[95], r3c[29], r3s[30], r3c[30]);

HA	inst1118	(r3s[1], pp[128], m[4], r4c[0]);
FA	inst1119	(r3s[2], pp[129], r4c[0], r4s[1], r4c[1]);
FA	inst1120	(r3s[3], pp[130], r4c[1], r4s[2], r4c[2]);
FA	inst1121	(r3s[4], pp[131], r4c[2], r4s[3], r4c[3]);
FA	inst1122	(r3s[5], pp[132], r4c[3], r4s[4], r4c[4]);
FA	inst1123	(r3s[6], pp[133], r4c[4], r4s[5], r4c[5]);
FA	inst1124	(r3s[7], pp[134], r4c[5], r4s[6], r4c[6]);
FA	inst1125	(r3s[8], pp[135], r4c[6], r4s[7], r4c[7]);
FA	inst1126	(r3s[9], pp[136], r4c[7], r4s[8], r4c[8]);
FA	inst1127	(r3s[10], pp[137], r4c[8], r4s[9], r4c[9]);
FA	inst1128	(r3s[11], pp[138], r4c[9], r4s[10], r4c[10]);
FA	inst1129	(r3s[12], pp[139], r4c[10], r4s[11], r4c[11]);
FA	inst1130	(r3s[13], pp[140], r4c[11], r4s[12], r4c[12]);
FA	inst1131	(r3s[14], pp[141], r4c[12], r4s[13], r4c[13]);
FA	inst1132	(r3s[15], pp[142], r4c[13], r4s[14], r4c[14]);
FA	inst1133	(r3s[16], pp[143], r4c[14], r4s[15], r4c[15]);
FA	inst1134	(r3s[17], pp[144], r4c[15], r4s[16], r4c[16]);
FA	inst1135	(r3s[18], pp[145], r4c[16], r4s[17], r4c[17]);
FA	inst1136	(r3s[19], pp[146], r4c[17], r4s[18], r4c[18]);
FA	inst1137	(r3s[20], pp[147], r4c[18], r4s[19], r4c[19]);
FA	inst1138	(r3s[21], pp[148], r4c[19], r4s[20], r4c[20]);
FA	inst1139	(r3s[22], pp[149], r4c[20], r4s[21], r4c[21]);
FA	inst1140	(r3s[23], pp[150], r4c[21], r4s[22], r4c[22]);
FA	inst1141	(r3s[24], pp[151], r4c[22], r4s[23], r4c[23]);
FA	inst1142	(r3s[25], pp[152], r4c[23], r4s[24], r4c[24]);
FA	inst1143	(r3s[26], pp[153], r4c[24], r4s[25], r4c[25]);
FA	inst1144	(r3s[27], pp[154], r4c[25], r4s[26], r4c[26]);
FA	inst1145	(r3s[28], pp[155], r4c[26], r4s[27], r4c[27]);
FA	inst1146	(r3s[29], pp[125], r4c[27], r4s[28], r4c[28]);
FA	inst1147	(r3s[30], pp[126], r4c[28], r4s[29], r4c[29]);
FA	inst1148	(r3c[30], pp[127], r4c[29], r4s[30], r4c[30]);

HA	inst1149	(r4s[1], pp[160], m[5], r5c[0]);
FA	inst1150	(r4s[2], pp[161], r5c[0], r5s[1], r5c[1]);
FA	inst1151	(r4s[3], pp[162], r5c[1], r5s[2], r5c[2]);
FA	inst1152	(r4s[4], pp[163], r5c[2], r5s[3], r5c[3]);
FA	inst1153	(r4s[5], pp[164], r5c[3], r5s[4], r5c[4]);
FA	inst1154	(r4s[6], pp[165], r5c[4], r5s[5], r5c[5]);
FA	inst1155	(r4s[7], pp[166], r5c[5], r5s[6], r5c[6]);
FA	inst1156	(r4s[8], pp[167], r5c[6], r5s[7], r5c[7]);
FA	inst1157	(r4s[9], pp[168], r5c[7], r5s[8], r5c[8]);
FA	inst1158	(r4s[10], pp[169], r5c[8], r5s[9], r5c[9]);
FA	inst1159	(r4s[11], pp[170], r5c[9], r5s[10], r5c[10]);
FA	inst1160	(r4s[12], pp[171], r5c[10], r5s[11], r5c[11]);
FA	inst1161	(r4s[13], pp[172], r5c[11], r5s[12], r5c[12]);
FA	inst1162	(r4s[14], pp[173], r5c[12], r5s[13], r5c[13]);
FA	inst1163	(r4s[15], pp[174], r5c[13], r5s[14], r5c[14]);
FA	inst1164	(r4s[16], pp[175], r5c[14], r5s[15], r5c[15]);
FA	inst1165	(r4s[17], pp[176], r5c[15], r5s[16], r5c[16]);
FA	inst1166	(r4s[18], pp[177], r5c[16], r5s[17], r5c[17]);
FA	inst1167	(r4s[19], pp[178], r5c[17], r5s[18], r5c[18]);
FA	inst1168	(r4s[20], pp[179], r5c[18], r5s[19], r5c[19]);
FA	inst1169	(r4s[21], pp[180], r5c[19], r5s[20], r5c[20]);
FA	inst1170	(r4s[22], pp[181], r5c[20], r5s[21], r5c[21]);
FA	inst1171	(r4s[23], pp[182], r5c[21], r5s[22], r5c[22]);
FA	inst1172	(r4s[24], pp[183], r5c[22], r5s[23], r5c[23]);
FA	inst1173	(r4s[25], pp[184], r5c[23], r5s[24], r5c[24]);
FA	inst1174	(r4s[26], pp[185], r5c[24], r5s[25], r5c[25]);
FA	inst1175	(r4s[27], pp[186], r5c[25], r5s[26], r5c[26]);
FA	inst1176	(r4s[28], pp[156], r5c[26], r5s[27], r5c[27]);
FA	inst1177	(r4s[29], pp[157], r5c[27], r5s[28], r5c[28]);
FA	inst1178	(r4s[30], pp[158], r5c[28], r5s[29], r5c[29]);
FA	inst1179	(r4c[30], pp[159], r5c[29], r5s[30], r5c[30]);

HA	inst1180	(r5s[1], pp[192], m[6], r6c[0]);
FA	inst1181	(r5s[2], pp[193], r6c[0], r6s[1], r6c[1]);
FA	inst1182	(r5s[3], pp[194], r6c[1], r6s[2], r6c[2]);
FA	inst1183	(r5s[4], pp[195], r6c[2], r6s[3], r6c[3]);
FA	inst1184	(r5s[5], pp[196], r6c[3], r6s[4], r6c[4]);
FA	inst1185	(r5s[6], pp[197], r6c[4], r6s[5], r6c[5]);
FA	inst1186	(r5s[7], pp[198], r6c[5], r6s[6], r6c[6]);
FA	inst1187	(r5s[8], pp[199], r6c[6], r6s[7], r6c[7]);
FA	inst1188	(r5s[9], pp[200], r6c[7], r6s[8], r6c[8]);
FA	inst1189	(r5s[10], pp[201], r6c[8], r6s[9], r6c[9]);
FA	inst1190	(r5s[11], pp[202], r6c[9], r6s[10], r6c[10]);
FA	inst1191	(r5s[12], pp[203], r6c[10], r6s[11], r6c[11]);
FA	inst1192	(r5s[13], pp[204], r6c[11], r6s[12], r6c[12]);
FA	inst1193	(r5s[14], pp[205], r6c[12], r6s[13], r6c[13]);
FA	inst1194	(r5s[15], pp[206], r6c[13], r6s[14], r6c[14]);
FA	inst1195	(r5s[16], pp[207], r6c[14], r6s[15], r6c[15]);
FA	inst1196	(r5s[17], pp[208], r6c[15], r6s[16], r6c[16]);
FA	inst1197	(r5s[18], pp[209], r6c[16], r6s[17], r6c[17]);
FA	inst1198	(r5s[19], pp[210], r6c[17], r6s[18], r6c[18]);
FA	inst1199	(r5s[20], pp[211], r6c[18], r6s[19], r6c[19]);
FA	inst1200	(r5s[21], pp[212], r6c[19], r6s[20], r6c[20]);
FA	inst1201	(r5s[22], pp[213], r6c[20], r6s[21], r6c[21]);
FA	inst1202	(r5s[23], pp[214], r6c[21], r6s[22], r6c[22]);
FA	inst1203	(r5s[24], pp[215], r6c[22], r6s[23], r6c[23]);
FA	inst1204	(r5s[25], pp[216], r6c[23], r6s[24], r6c[24]);
FA	inst1205	(r5s[26], pp[217], r6c[24], r6s[25], r6c[25]);
FA	inst1206	(r5s[27], pp[187], r6c[25], r6s[26], r6c[26]);
FA	inst1207	(r5s[28], pp[188], r6c[26], r6s[27], r6c[27]);
FA	inst1208	(r5s[29], pp[189], r6c[27], r6s[28], r6c[28]);
FA	inst1209	(r5s[30], pp[190], r6c[28], r6s[29], r6c[29]);
FA	inst1210	(r5c[30], pp[191], r6c[29], r6s[30], r6c[30]);

HA	inst1211	(r6s[1], pp[224], m[7], r7c[0]);
FA	inst1212	(r6s[2], pp[225], r7c[0], r7s[1], r7c[1]);
FA	inst1213	(r6s[3], pp[226], r7c[1], r7s[2], r7c[2]);
FA	inst1214	(r6s[4], pp[227], r7c[2], r7s[3], r7c[3]);
FA	inst1215	(r6s[5], pp[228], r7c[3], r7s[4], r7c[4]);
FA	inst1216	(r6s[6], pp[229], r7c[4], r7s[5], r7c[5]);
FA	inst1217	(r6s[7], pp[230], r7c[5], r7s[6], r7c[6]);
FA	inst1218	(r6s[8], pp[231], r7c[6], r7s[7], r7c[7]);
FA	inst1219	(r6s[9], pp[232], r7c[7], r7s[8], r7c[8]);
FA	inst1220	(r6s[10], pp[233], r7c[8], r7s[9], r7c[9]);
FA	inst1221	(r6s[11], pp[234], r7c[9], r7s[10], r7c[10]);
FA	inst1222	(r6s[12], pp[235], r7c[10], r7s[11], r7c[11]);
FA	inst1223	(r6s[13], pp[236], r7c[11], r7s[12], r7c[12]);
FA	inst1224	(r6s[14], pp[237], r7c[12], r7s[13], r7c[13]);
FA	inst1225	(r6s[15], pp[238], r7c[13], r7s[14], r7c[14]);
FA	inst1226	(r6s[16], pp[239], r7c[14], r7s[15], r7c[15]);
FA	inst1227	(r6s[17], pp[240], r7c[15], r7s[16], r7c[16]);
FA	inst1228	(r6s[18], pp[241], r7c[16], r7s[17], r7c[17]);
FA	inst1229	(r6s[19], pp[242], r7c[17], r7s[18], r7c[18]);
FA	inst1230	(r6s[20], pp[243], r7c[18], r7s[19], r7c[19]);
FA	inst1231	(r6s[21], pp[244], r7c[19], r7s[20], r7c[20]);
FA	inst1232	(r6s[22], pp[245], r7c[20], r7s[21], r7c[21]);
FA	inst1233	(r6s[23], pp[246], r7c[21], r7s[22], r7c[22]);
FA	inst1234	(r6s[24], pp[247], r7c[22], r7s[23], r7c[23]);
FA	inst1235	(r6s[25], pp[248], r7c[23], r7s[24], r7c[24]);
FA	inst1236	(r6s[26], pp[218], r7c[24], r7s[25], r7c[25]);
FA	inst1237	(r6s[27], pp[219], r7c[25], r7s[26], r7c[26]);
FA	inst1238	(r6s[28], pp[220], r7c[26], r7s[27], r7c[27]);
FA	inst1239	(r6s[29], pp[221], r7c[27], r7s[28], r7c[28]);
FA	inst1240	(r6s[30], pp[222], r7c[28], r7s[29], r7c[29]);
FA	inst1241	(r6c[30], pp[223], r7c[29], r7s[30], r7c[30]);

HA	inst1242	(r7s[1], pp[256], m[8], r8c[0]);
FA	inst1243	(r7s[2], pp[257], r8c[0], r8s[1], r8c[1]);
FA	inst1244	(r7s[3], pp[258], r8c[1], r8s[2], r8c[2]);
FA	inst1245	(r7s[4], pp[259], r8c[2], r8s[3], r8c[3]);
FA	inst1246	(r7s[5], pp[260], r8c[3], r8s[4], r8c[4]);
FA	inst1247	(r7s[6], pp[261], r8c[4], r8s[5], r8c[5]);
FA	inst1248	(r7s[7], pp[262], r8c[5], r8s[6], r8c[6]);
FA	inst1249	(r7s[8], pp[263], r8c[6], r8s[7], r8c[7]);
FA	inst1250	(r7s[9], pp[264], r8c[7], r8s[8], r8c[8]);
FA	inst1251	(r7s[10], pp[265], r8c[8], r8s[9], r8c[9]);
FA	inst1252	(r7s[11], pp[266], r8c[9], r8s[10], r8c[10]);
FA	inst1253	(r7s[12], pp[267], r8c[10], r8s[11], r8c[11]);
FA	inst1254	(r7s[13], pp[268], r8c[11], r8s[12], r8c[12]);
FA	inst1255	(r7s[14], pp[269], r8c[12], r8s[13], r8c[13]);
FA	inst1256	(r7s[15], pp[270], r8c[13], r8s[14], r8c[14]);
FA	inst1257	(r7s[16], pp[271], r8c[14], r8s[15], r8c[15]);
FA	inst1258	(r7s[17], pp[272], r8c[15], r8s[16], r8c[16]);
FA	inst1259	(r7s[18], pp[273], r8c[16], r8s[17], r8c[17]);
FA	inst1260	(r7s[19], pp[274], r8c[17], r8s[18], r8c[18]);
FA	inst1261	(r7s[20], pp[275], r8c[18], r8s[19], r8c[19]);
FA	inst1262	(r7s[21], pp[276], r8c[19], r8s[20], r8c[20]);
FA	inst1263	(r7s[22], pp[277], r8c[20], r8s[21], r8c[21]);
FA	inst1264	(r7s[23], pp[278], r8c[21], r8s[22], r8c[22]);
FA	inst1265	(r7s[24], pp[279], r8c[22], r8s[23], r8c[23]);
FA	inst1266	(r7s[25], pp[249], r8c[23], r8s[24], r8c[24]);
FA	inst1267	(r7s[26], pp[250], r8c[24], r8s[25], r8c[25]);
FA	inst1268	(r7s[27], pp[251], r8c[25], r8s[26], r8c[26]);
FA	inst1269	(r7s[28], pp[252], r8c[26], r8s[27], r8c[27]);
FA	inst1270	(r7s[29], pp[253], r8c[27], r8s[28], r8c[28]);
FA	inst1271	(r7s[30], pp[254], r8c[28], r8s[29], r8c[29]);
FA	inst1272	(r7c[30], pp[255], r8c[29], r8s[30], r8c[30]);

HA	inst1273	(r8s[1], pp[288], m[9], r9c[0]);
FA	inst1274	(r8s[2], pp[289], r9c[0], r9s[1], r9c[1]);
FA	inst1275	(r8s[3], pp[290], r9c[1], r9s[2], r9c[2]);
FA	inst1276	(r8s[4], pp[291], r9c[2], r9s[3], r9c[3]);
FA	inst1277	(r8s[5], pp[292], r9c[3], r9s[4], r9c[4]);
FA	inst1278	(r8s[6], pp[293], r9c[4], r9s[5], r9c[5]);
FA	inst1279	(r8s[7], pp[294], r9c[5], r9s[6], r9c[6]);
FA	inst1280	(r8s[8], pp[295], r9c[6], r9s[7], r9c[7]);
FA	inst1281	(r8s[9], pp[296], r9c[7], r9s[8], r9c[8]);
FA	inst1282	(r8s[10], pp[297], r9c[8], r9s[9], r9c[9]);
FA	inst1283	(r8s[11], pp[298], r9c[9], r9s[10], r9c[10]);
FA	inst1284	(r8s[12], pp[299], r9c[10], r9s[11], r9c[11]);
FA	inst1285	(r8s[13], pp[300], r9c[11], r9s[12], r9c[12]);
FA	inst1286	(r8s[14], pp[301], r9c[12], r9s[13], r9c[13]);
FA	inst1287	(r8s[15], pp[302], r9c[13], r9s[14], r9c[14]);
FA	inst1288	(r8s[16], pp[303], r9c[14], r9s[15], r9c[15]);
FA	inst1289	(r8s[17], pp[304], r9c[15], r9s[16], r9c[16]);
FA	inst1290	(r8s[18], pp[305], r9c[16], r9s[17], r9c[17]);
FA	inst1291	(r8s[19], pp[306], r9c[17], r9s[18], r9c[18]);
FA	inst1292	(r8s[20], pp[307], r9c[18], r9s[19], r9c[19]);
FA	inst1293	(r8s[21], pp[308], r9c[19], r9s[20], r9c[20]);
FA	inst1294	(r8s[22], pp[309], r9c[20], r9s[21], r9c[21]);
FA	inst1295	(r8s[23], pp[310], r9c[21], r9s[22], r9c[22]);
FA	inst1296	(r8s[24], pp[280], r9c[22], r9s[23], r9c[23]);
FA	inst1297	(r8s[25], pp[281], r9c[23], r9s[24], r9c[24]);
FA	inst1298	(r8s[26], pp[282], r9c[24], r9s[25], r9c[25]);
FA	inst1299	(r8s[27], pp[283], r9c[25], r9s[26], r9c[26]);
FA	inst1300	(r8s[28], pp[284], r9c[26], r9s[27], r9c[27]);
FA	inst1301	(r8s[29], pp[285], r9c[27], r9s[28], r9c[28]);
FA	inst1302	(r8s[30], pp[286], r9c[28], r9s[29], r9c[29]);
FA	inst1303	(r8c[30], pp[287], r9c[29], r9s[30], r9c[30]);

HA	inst1304	(r9s[1], pp[320], m[10], r10c[0]);
FA	inst1305	(r9s[2], pp[321], r10c[0], r10s[1], r10c[1]);
FA	inst1306	(r9s[3], pp[322], r10c[1], r10s[2], r10c[2]);
FA	inst1307	(r9s[4], pp[323], r10c[2], r10s[3], r10c[3]);
FA	inst1308	(r9s[5], pp[324], r10c[3], r10s[4], r10c[4]);
FA	inst1309	(r9s[6], pp[325], r10c[4], r10s[5], r10c[5]);
FA	inst1310	(r9s[7], pp[326], r10c[5], r10s[6], r10c[6]);
FA	inst1311	(r9s[8], pp[327], r10c[6], r10s[7], r10c[7]);
FA	inst1312	(r9s[9], pp[328], r10c[7], r10s[8], r10c[8]);
FA	inst1313	(r9s[10], pp[329], r10c[8], r10s[9], r10c[9]);
FA	inst1314	(r9s[11], pp[330], r10c[9], r10s[10], r10c[10]);
FA	inst1315	(r9s[12], pp[331], r10c[10], r10s[11], r10c[11]);
FA	inst1316	(r9s[13], pp[332], r10c[11], r10s[12], r10c[12]);
FA	inst1317	(r9s[14], pp[333], r10c[12], r10s[13], r10c[13]);
FA	inst1318	(r9s[15], pp[334], r10c[13], r10s[14], r10c[14]);
FA	inst1319	(r9s[16], pp[335], r10c[14], r10s[15], r10c[15]);
FA	inst1320	(r9s[17], pp[336], r10c[15], r10s[16], r10c[16]);
FA	inst1321	(r9s[18], pp[337], r10c[16], r10s[17], r10c[17]);
FA	inst1322	(r9s[19], pp[338], r10c[17], r10s[18], r10c[18]);
FA	inst1323	(r9s[20], pp[339], r10c[18], r10s[19], r10c[19]);
FA	inst1324	(r9s[21], pp[340], r10c[19], r10s[20], r10c[20]);
FA	inst1325	(r9s[22], pp[341], r10c[20], r10s[21], r10c[21]);
FA	inst1326	(r9s[23], pp[311], r10c[21], r10s[22], r10c[22]);
FA	inst1327	(r9s[24], pp[312], r10c[22], r10s[23], r10c[23]);
FA	inst1328	(r9s[25], pp[313], r10c[23], r10s[24], r10c[24]);
FA	inst1329	(r9s[26], pp[314], r10c[24], r10s[25], r10c[25]);
FA	inst1330	(r9s[27], pp[315], r10c[25], r10s[26], r10c[26]);
FA	inst1331	(r9s[28], pp[316], r10c[26], r10s[27], r10c[27]);
FA	inst1332	(r9s[29], pp[317], r10c[27], r10s[28], r10c[28]);
FA	inst1333	(r9s[30], pp[318], r10c[28], r10s[29], r10c[29]);
FA	inst1334	(r9c[30], pp[319], r10c[29], r10s[30], r10c[30]);

HA	inst1335	(r10s[1], pp[352], m[11], r11c[0]);
FA	inst1336	(r10s[2], pp[353], r11c[0], r11s[1], r11c[1]);
FA	inst1337	(r10s[3], pp[354], r11c[1], r11s[2], r11c[2]);
FA	inst1338	(r10s[4], pp[355], r11c[2], r11s[3], r11c[3]);
FA	inst1339	(r10s[5], pp[356], r11c[3], r11s[4], r11c[4]);
FA	inst1340	(r10s[6], pp[357], r11c[4], r11s[5], r11c[5]);
FA	inst1341	(r10s[7], pp[358], r11c[5], r11s[6], r11c[6]);
FA	inst1342	(r10s[8], pp[359], r11c[6], r11s[7], r11c[7]);
FA	inst1343	(r10s[9], pp[360], r11c[7], r11s[8], r11c[8]);
FA	inst1344	(r10s[10], pp[361], r11c[8], r11s[9], r11c[9]);
FA	inst1345	(r10s[11], pp[362], r11c[9], r11s[10], r11c[10]);
FA	inst1346	(r10s[12], pp[363], r11c[10], r11s[11], r11c[11]);
FA	inst1347	(r10s[13], pp[364], r11c[11], r11s[12], r11c[12]);
FA	inst1348	(r10s[14], pp[365], r11c[12], r11s[13], r11c[13]);
FA	inst1349	(r10s[15], pp[366], r11c[13], r11s[14], r11c[14]);
FA	inst1350	(r10s[16], pp[367], r11c[14], r11s[15], r11c[15]);
FA	inst1351	(r10s[17], pp[368], r11c[15], r11s[16], r11c[16]);
FA	inst1352	(r10s[18], pp[369], r11c[16], r11s[17], r11c[17]);
FA	inst1353	(r10s[19], pp[370], r11c[17], r11s[18], r11c[18]);
FA	inst1354	(r10s[20], pp[371], r11c[18], r11s[19], r11c[19]);
FA	inst1355	(r10s[21], pp[372], r11c[19], r11s[20], r11c[20]);
FA	inst1356	(r10s[22], pp[342], r11c[20], r11s[21], r11c[21]);
FA	inst1357	(r10s[23], pp[343], r11c[21], r11s[22], r11c[22]);
FA	inst1358	(r10s[24], pp[344], r11c[22], r11s[23], r11c[23]);
FA	inst1359	(r10s[25], pp[345], r11c[23], r11s[24], r11c[24]);
FA	inst1360	(r10s[26], pp[346], r11c[24], r11s[25], r11c[25]);
FA	inst1361	(r10s[27], pp[347], r11c[25], r11s[26], r11c[26]);
FA	inst1362	(r10s[28], pp[348], r11c[26], r11s[27], r11c[27]);
FA	inst1363	(r10s[29], pp[349], r11c[27], r11s[28], r11c[28]);
FA	inst1364	(r10s[30], pp[350], r11c[28], r11s[29], r11c[29]);
FA	inst1365	(r10c[30], pp[351], r11c[29], r11s[30], r11c[30]);

HA	inst1366	(r11s[1], pp[384], m[12], r12c[0]);
FA	inst1367	(r11s[2], pp[385], r12c[0], r12s[1], r12c[1]);
FA	inst1368	(r11s[3], pp[386], r12c[1], r12s[2], r12c[2]);
FA	inst1369	(r11s[4], pp[387], r12c[2], r12s[3], r12c[3]);
FA	inst1370	(r11s[5], pp[388], r12c[3], r12s[4], r12c[4]);
FA	inst1371	(r11s[6], pp[389], r12c[4], r12s[5], r12c[5]);
FA	inst1372	(r11s[7], pp[390], r12c[5], r12s[6], r12c[6]);
FA	inst1373	(r11s[8], pp[391], r12c[6], r12s[7], r12c[7]);
FA	inst1374	(r11s[9], pp[392], r12c[7], r12s[8], r12c[8]);
FA	inst1375	(r11s[10], pp[393], r12c[8], r12s[9], r12c[9]);
FA	inst1376	(r11s[11], pp[394], r12c[9], r12s[10], r12c[10]);
FA	inst1377	(r11s[12], pp[395], r12c[10], r12s[11], r12c[11]);
FA	inst1378	(r11s[13], pp[396], r12c[11], r12s[12], r12c[12]);
FA	inst1379	(r11s[14], pp[397], r12c[12], r12s[13], r12c[13]);
FA	inst1380	(r11s[15], pp[398], r12c[13], r12s[14], r12c[14]);
FA	inst1381	(r11s[16], pp[399], r12c[14], r12s[15], r12c[15]);
FA	inst1382	(r11s[17], pp[400], r12c[15], r12s[16], r12c[16]);
FA	inst1383	(r11s[18], pp[401], r12c[16], r12s[17], r12c[17]);
FA	inst1384	(r11s[19], pp[402], r12c[17], r12s[18], r12c[18]);
FA	inst1385	(r11s[20], pp[403], r12c[18], r12s[19], r12c[19]);
FA	inst1386	(r11s[21], pp[373], r12c[19], r12s[20], r12c[20]);
FA	inst1387	(r11s[22], pp[374], r12c[20], r12s[21], r12c[21]);
FA	inst1388	(r11s[23], pp[375], r12c[21], r12s[22], r12c[22]);
FA	inst1389	(r11s[24], pp[376], r12c[22], r12s[23], r12c[23]);
FA	inst1390	(r11s[25], pp[377], r12c[23], r12s[24], r12c[24]);
FA	inst1391	(r11s[26], pp[378], r12c[24], r12s[25], r12c[25]);
FA	inst1392	(r11s[27], pp[379], r12c[25], r12s[26], r12c[26]);
FA	inst1393	(r11s[28], pp[380], r12c[26], r12s[27], r12c[27]);
FA	inst1394	(r11s[29], pp[381], r12c[27], r12s[28], r12c[28]);
FA	inst1395	(r11s[30], pp[382], r12c[28], r12s[29], r12c[29]);
FA	inst1396	(r11c[30], pp[383], r12c[29], r12s[30], r12c[30]);

HA	inst1397	(r12s[1], pp[416], m[13], r13c[0]);
FA	inst1398	(r12s[2], pp[417], r13c[0], r13s[1], r13c[1]);
FA	inst1399	(r12s[3], pp[418], r13c[1], r13s[2], r13c[2]);
FA	inst1400	(r12s[4], pp[419], r13c[2], r13s[3], r13c[3]);
FA	inst1401	(r12s[5], pp[420], r13c[3], r13s[4], r13c[4]);
FA	inst1402	(r12s[6], pp[421], r13c[4], r13s[5], r13c[5]);
FA	inst1403	(r12s[7], pp[422], r13c[5], r13s[6], r13c[6]);
FA	inst1404	(r12s[8], pp[423], r13c[6], r13s[7], r13c[7]);
FA	inst1405	(r12s[9], pp[424], r13c[7], r13s[8], r13c[8]);
FA	inst1406	(r12s[10], pp[425], r13c[8], r13s[9], r13c[9]);
FA	inst1407	(r12s[11], pp[426], r13c[9], r13s[10], r13c[10]);
FA	inst1408	(r12s[12], pp[427], r13c[10], r13s[11], r13c[11]);
FA	inst1409	(r12s[13], pp[428], r13c[11], r13s[12], r13c[12]);
FA	inst1410	(r12s[14], pp[429], r13c[12], r13s[13], r13c[13]);
FA	inst1411	(r12s[15], pp[430], r13c[13], r13s[14], r13c[14]);
FA	inst1412	(r12s[16], pp[431], r13c[14], r13s[15], r13c[15]);
FA	inst1413	(r12s[17], pp[432], r13c[15], r13s[16], r13c[16]);
FA	inst1414	(r12s[18], pp[433], r13c[16], r13s[17], r13c[17]);
FA	inst1415	(r12s[19], pp[434], r13c[17], r13s[18], r13c[18]);
FA	inst1416	(r12s[20], pp[404], r13c[18], r13s[19], r13c[19]);
FA	inst1417	(r12s[21], pp[405], r13c[19], r13s[20], r13c[20]);
FA	inst1418	(r12s[22], pp[406], r13c[20], r13s[21], r13c[21]);
FA	inst1419	(r12s[23], pp[407], r13c[21], r13s[22], r13c[22]);
FA	inst1420	(r12s[24], pp[408], r13c[22], r13s[23], r13c[23]);
FA	inst1421	(r12s[25], pp[409], r13c[23], r13s[24], r13c[24]);
FA	inst1422	(r12s[26], pp[410], r13c[24], r13s[25], r13c[25]);
FA	inst1423	(r12s[27], pp[411], r13c[25], r13s[26], r13c[26]);
FA	inst1424	(r12s[28], pp[412], r13c[26], r13s[27], r13c[27]);
FA	inst1425	(r12s[29], pp[413], r13c[27], r13s[28], r13c[28]);
FA	inst1426	(r12s[30], pp[414], r13c[28], r13s[29], r13c[29]);
FA	inst1427	(r12c[30], pp[415], r13c[29], r13s[30], r13c[30]);

HA	inst1428	(r13s[1], pp[448], m[14], r14c[0]);
FA	inst1429	(r13s[2], pp[449], r14c[0], r14s[1], r14c[1]);
FA	inst1430	(r13s[3], pp[450], r14c[1], r14s[2], r14c[2]);
FA	inst1431	(r13s[4], pp[451], r14c[2], r14s[3], r14c[3]);
FA	inst1432	(r13s[5], pp[452], r14c[3], r14s[4], r14c[4]);
FA	inst1433	(r13s[6], pp[453], r14c[4], r14s[5], r14c[5]);
FA	inst1434	(r13s[7], pp[454], r14c[5], r14s[6], r14c[6]);
FA	inst1435	(r13s[8], pp[455], r14c[6], r14s[7], r14c[7]);
FA	inst1436	(r13s[9], pp[456], r14c[7], r14s[8], r14c[8]);
FA	inst1437	(r13s[10], pp[457], r14c[8], r14s[9], r14c[9]);
FA	inst1438	(r13s[11], pp[458], r14c[9], r14s[10], r14c[10]);
FA	inst1439	(r13s[12], pp[459], r14c[10], r14s[11], r14c[11]);
FA	inst1440	(r13s[13], pp[460], r14c[11], r14s[12], r14c[12]);
FA	inst1441	(r13s[14], pp[461], r14c[12], r14s[13], r14c[13]);
FA	inst1442	(r13s[15], pp[462], r14c[13], r14s[14], r14c[14]);
FA	inst1443	(r13s[16], pp[463], r14c[14], r14s[15], r14c[15]);
FA	inst1444	(r13s[17], pp[464], r14c[15], r14s[16], r14c[16]);
FA	inst1445	(r13s[18], pp[465], r14c[16], r14s[17], r14c[17]);
FA	inst1446	(r13s[19], pp[435], r14c[17], r14s[18], r14c[18]);
FA	inst1447	(r13s[20], pp[436], r14c[18], r14s[19], r14c[19]);
FA	inst1448	(r13s[21], pp[437], r14c[19], r14s[20], r14c[20]);
FA	inst1449	(r13s[22], pp[438], r14c[20], r14s[21], r14c[21]);
FA	inst1450	(r13s[23], pp[439], r14c[21], r14s[22], r14c[22]);
FA	inst1451	(r13s[24], pp[440], r14c[22], r14s[23], r14c[23]);
FA	inst1452	(r13s[25], pp[441], r14c[23], r14s[24], r14c[24]);
FA	inst1453	(r13s[26], pp[442], r14c[24], r14s[25], r14c[25]);
FA	inst1454	(r13s[27], pp[443], r14c[25], r14s[26], r14c[26]);
FA	inst1455	(r13s[28], pp[444], r14c[26], r14s[27], r14c[27]);
FA	inst1456	(r13s[29], pp[445], r14c[27], r14s[28], r14c[28]);
FA	inst1457	(r13s[30], pp[446], r14c[28], r14s[29], r14c[29]);
FA	inst1458	(r13c[30], pp[447], r14c[29], r14s[30], r14c[30]);

HA	inst1459	(r14s[1], pp[480], m[15], r15c[0]);
FA	inst1460	(r14s[2], pp[481], r15c[0], r15s[1], r15c[1]);
FA	inst1461	(r14s[3], pp[482], r15c[1], r15s[2], r15c[2]);
FA	inst1462	(r14s[4], pp[483], r15c[2], r15s[3], r15c[3]);
FA	inst1463	(r14s[5], pp[484], r15c[3], r15s[4], r15c[4]);
FA	inst1464	(r14s[6], pp[485], r15c[4], r15s[5], r15c[5]);
FA	inst1465	(r14s[7], pp[486], r15c[5], r15s[6], r15c[6]);
FA	inst1466	(r14s[8], pp[487], r15c[6], r15s[7], r15c[7]);
FA	inst1467	(r14s[9], pp[488], r15c[7], r15s[8], r15c[8]);
FA	inst1468	(r14s[10], pp[489], r15c[8], r15s[9], r15c[9]);
FA	inst1469	(r14s[11], pp[490], r15c[9], r15s[10], r15c[10]);
FA	inst1470	(r14s[12], pp[491], r15c[10], r15s[11], r15c[11]);
FA	inst1471	(r14s[13], pp[492], r15c[11], r15s[12], r15c[12]);
FA	inst1472	(r14s[14], pp[493], r15c[12], r15s[13], r15c[13]);
FA	inst1473	(r14s[15], pp[494], r15c[13], r15s[14], r15c[14]);
FA	inst1474	(r14s[16], pp[495], r15c[14], r15s[15], r15c[15]);
FA	inst1475	(r14s[17], pp[496], r15c[15], r15s[16], r15c[16]);
FA	inst1476	(r14s[18], pp[466], r15c[16], r15s[17], r15c[17]);
FA	inst1477	(r14s[19], pp[467], r15c[17], r15s[18], r15c[18]);
FA	inst1478	(r14s[20], pp[468], r15c[18], r15s[19], r15c[19]);
FA	inst1479	(r14s[21], pp[469], r15c[19], r15s[20], r15c[20]);
FA	inst1480	(r14s[22], pp[470], r15c[20], r15s[21], r15c[21]);
FA	inst1481	(r14s[23], pp[471], r15c[21], r15s[22], r15c[22]);
FA	inst1482	(r14s[24], pp[472], r15c[22], r15s[23], r15c[23]);
FA	inst1483	(r14s[25], pp[473], r15c[23], r15s[24], r15c[24]);
FA	inst1484	(r14s[26], pp[474], r15c[24], r15s[25], r15c[25]);
FA	inst1485	(r14s[27], pp[475], r15c[25], r15s[26], r15c[26]);
FA	inst1486	(r14s[28], pp[476], r15c[26], r15s[27], r15c[27]);
FA	inst1487	(r14s[29], pp[477], r15c[27], r15s[28], r15c[28]);
FA	inst1488	(r14s[30], pp[478], r15c[28], r15s[29], r15c[29]);
FA	inst1489	(r14c[30], pp[479], r15c[29], r15s[30], r15c[30]);

HA	inst1490	(r15s[1], pp[512], m[16], r16c[0]);
FA	inst1491	(r15s[2], pp[513], r16c[0], r16s[1], r16c[1]);
FA	inst1492	(r15s[3], pp[514], r16c[1], r16s[2], r16c[2]);
FA	inst1493	(r15s[4], pp[515], r16c[2], r16s[3], r16c[3]);
FA	inst1494	(r15s[5], pp[516], r16c[3], r16s[4], r16c[4]);
FA	inst1495	(r15s[6], pp[517], r16c[4], r16s[5], r16c[5]);
FA	inst1496	(r15s[7], pp[518], r16c[5], r16s[6], r16c[6]);
FA	inst1497	(r15s[8], pp[519], r16c[6], r16s[7], r16c[7]);
FA	inst1498	(r15s[9], pp[520], r16c[7], r16s[8], r16c[8]);
FA	inst1499	(r15s[10], pp[521], r16c[8], r16s[9], r16c[9]);
FA	inst1500	(r15s[11], pp[522], r16c[9], r16s[10], r16c[10]);
FA	inst1501	(r15s[12], pp[523], r16c[10], r16s[11], r16c[11]);
FA	inst1502	(r15s[13], pp[524], r16c[11], r16s[12], r16c[12]);
FA	inst1503	(r15s[14], pp[525], r16c[12], r16s[13], r16c[13]);
FA	inst1504	(r15s[15], pp[526], r16c[13], r16s[14], r16c[14]);
FA	inst1505	(r15s[16], pp[527], r16c[14], r16s[15], r16c[15]);
FA	inst1506	(r15s[17], pp[497], r16c[15], r16s[16], r16c[16]);
FA	inst1507	(r15s[18], pp[498], r16c[16], r16s[17], r16c[17]);
FA	inst1508	(r15s[19], pp[499], r16c[17], r16s[18], r16c[18]);
FA	inst1509	(r15s[20], pp[500], r16c[18], r16s[19], r16c[19]);
FA	inst1510	(r15s[21], pp[501], r16c[19], r16s[20], r16c[20]);
FA	inst1511	(r15s[22], pp[502], r16c[20], r16s[21], r16c[21]);
FA	inst1512	(r15s[23], pp[503], r16c[21], r16s[22], r16c[22]);
FA	inst1513	(r15s[24], pp[504], r16c[22], r16s[23], r16c[23]);
FA	inst1514	(r15s[25], pp[505], r16c[23], r16s[24], r16c[24]);
FA	inst1515	(r15s[26], pp[506], r16c[24], r16s[25], r16c[25]);
FA	inst1516	(r15s[27], pp[507], r16c[25], r16s[26], r16c[26]);
FA	inst1517	(r15s[28], pp[508], r16c[26], r16s[27], r16c[27]);
FA	inst1518	(r15s[29], pp[509], r16c[27], r16s[28], r16c[28]);
FA	inst1519	(r15s[30], pp[510], r16c[28], r16s[29], r16c[29]);
FA	inst1520	(r15c[30], pp[511], r16c[29], r16s[30], r16c[30]);

HA	inst1521	(r16s[1], pp[544], m[17], r17c[0]);
FA	inst1522	(r16s[2], pp[545], r17c[0], r17s[1], r17c[1]);
FA	inst1523	(r16s[3], pp[546], r17c[1], r17s[2], r17c[2]);
FA	inst1524	(r16s[4], pp[547], r17c[2], r17s[3], r17c[3]);
FA	inst1525	(r16s[5], pp[548], r17c[3], r17s[4], r17c[4]);
FA	inst1526	(r16s[6], pp[549], r17c[4], r17s[5], r17c[5]);
FA	inst1527	(r16s[7], pp[550], r17c[5], r17s[6], r17c[6]);
FA	inst1528	(r16s[8], pp[551], r17c[6], r17s[7], r17c[7]);
FA	inst1529	(r16s[9], pp[552], r17c[7], r17s[8], r17c[8]);
FA	inst1530	(r16s[10], pp[553], r17c[8], r17s[9], r17c[9]);
FA	inst1531	(r16s[11], pp[554], r17c[9], r17s[10], r17c[10]);
FA	inst1532	(r16s[12], pp[555], r17c[10], r17s[11], r17c[11]);
FA	inst1533	(r16s[13], pp[556], r17c[11], r17s[12], r17c[12]);
FA	inst1534	(r16s[14], pp[557], r17c[12], r17s[13], r17c[13]);
FA	inst1535	(r16s[15], pp[558], r17c[13], r17s[14], r17c[14]);
FA	inst1536	(r16s[16], pp[528], r17c[14], r17s[15], r17c[15]);
FA	inst1537	(r16s[17], pp[529], r17c[15], r17s[16], r17c[16]);
FA	inst1538	(r16s[18], pp[530], r17c[16], r17s[17], r17c[17]);
FA	inst1539	(r16s[19], pp[531], r17c[17], r17s[18], r17c[18]);
FA	inst1540	(r16s[20], pp[532], r17c[18], r17s[19], r17c[19]);
FA	inst1541	(r16s[21], pp[533], r17c[19], r17s[20], r17c[20]);
FA	inst1542	(r16s[22], pp[534], r17c[20], r17s[21], r17c[21]);
FA	inst1543	(r16s[23], pp[535], r17c[21], r17s[22], r17c[22]);
FA	inst1544	(r16s[24], pp[536], r17c[22], r17s[23], r17c[23]);
FA	inst1545	(r16s[25], pp[537], r17c[23], r17s[24], r17c[24]);
FA	inst1546	(r16s[26], pp[538], r17c[24], r17s[25], r17c[25]);
FA	inst1547	(r16s[27], pp[539], r17c[25], r17s[26], r17c[26]);
FA	inst1548	(r16s[28], pp[540], r17c[26], r17s[27], r17c[27]);
FA	inst1549	(r16s[29], pp[541], r17c[27], r17s[28], r17c[28]);
FA	inst1550	(r16s[30], pp[542], r17c[28], r17s[29], r17c[29]);
FA	inst1551	(r16c[30], pp[543], r17c[29], r17s[30], r17c[30]);

HA	inst1552	(r17s[1], pp[576], m[18], r18c[0]);
FA	inst1553	(r17s[2], pp[577], r18c[0], r18s[1], r18c[1]);
FA	inst1554	(r17s[3], pp[578], r18c[1], r18s[2], r18c[2]);
FA	inst1555	(r17s[4], pp[579], r18c[2], r18s[3], r18c[3]);
FA	inst1556	(r17s[5], pp[580], r18c[3], r18s[4], r18c[4]);
FA	inst1557	(r17s[6], pp[581], r18c[4], r18s[5], r18c[5]);
FA	inst1558	(r17s[7], pp[582], r18c[5], r18s[6], r18c[6]);
FA	inst1559	(r17s[8], pp[583], r18c[6], r18s[7], r18c[7]);
FA	inst1560	(r17s[9], pp[584], r18c[7], r18s[8], r18c[8]);
FA	inst1561	(r17s[10], pp[585], r18c[8], r18s[9], r18c[9]);
FA	inst1562	(r17s[11], pp[586], r18c[9], r18s[10], r18c[10]);
FA	inst1563	(r17s[12], pp[587], r18c[10], r18s[11], r18c[11]);
FA	inst1564	(r17s[13], pp[588], r18c[11], r18s[12], r18c[12]);
FA	inst1565	(r17s[14], pp[589], r18c[12], r18s[13], r18c[13]);
FA	inst1566	(r17s[15], pp[559], r18c[13], r18s[14], r18c[14]);
FA	inst1567	(r17s[16], pp[560], r18c[14], r18s[15], r18c[15]);
FA	inst1568	(r17s[17], pp[561], r18c[15], r18s[16], r18c[16]);
FA	inst1569	(r17s[18], pp[562], r18c[16], r18s[17], r18c[17]);
FA	inst1570	(r17s[19], pp[563], r18c[17], r18s[18], r18c[18]);
FA	inst1571	(r17s[20], pp[564], r18c[18], r18s[19], r18c[19]);
FA	inst1572	(r17s[21], pp[565], r18c[19], r18s[20], r18c[20]);
FA	inst1573	(r17s[22], pp[566], r18c[20], r18s[21], r18c[21]);
FA	inst1574	(r17s[23], pp[567], r18c[21], r18s[22], r18c[22]);
FA	inst1575	(r17s[24], pp[568], r18c[22], r18s[23], r18c[23]);
FA	inst1576	(r17s[25], pp[569], r18c[23], r18s[24], r18c[24]);
FA	inst1577	(r17s[26], pp[570], r18c[24], r18s[25], r18c[25]);
FA	inst1578	(r17s[27], pp[571], r18c[25], r18s[26], r18c[26]);
FA	inst1579	(r17s[28], pp[572], r18c[26], r18s[27], r18c[27]);
FA	inst1580	(r17s[29], pp[573], r18c[27], r18s[28], r18c[28]);
FA	inst1581	(r17s[30], pp[574], r18c[28], r18s[29], r18c[29]);
FA	inst1582	(r17c[30], pp[575], r18c[29], r18s[30], r18c[30]);

HA	inst1583	(r18s[1], pp[608], m[19], r19c[0]);
FA	inst1584	(r18s[2], pp[609], r19c[0], r19s[1], r19c[1]);
FA	inst1585	(r18s[3], pp[610], r19c[1], r19s[2], r19c[2]);
FA	inst1586	(r18s[4], pp[611], r19c[2], r19s[3], r19c[3]);
FA	inst1587	(r18s[5], pp[612], r19c[3], r19s[4], r19c[4]);
FA	inst1588	(r18s[6], pp[613], r19c[4], r19s[5], r19c[5]);
FA	inst1589	(r18s[7], pp[614], r19c[5], r19s[6], r19c[6]);
FA	inst1590	(r18s[8], pp[615], r19c[6], r19s[7], r19c[7]);
FA	inst1591	(r18s[9], pp[616], r19c[7], r19s[8], r19c[8]);
FA	inst1592	(r18s[10], pp[617], r19c[8], r19s[9], r19c[9]);
FA	inst1593	(r18s[11], pp[618], r19c[9], r19s[10], r19c[10]);
FA	inst1594	(r18s[12], pp[619], r19c[10], r19s[11], r19c[11]);
FA	inst1595	(r18s[13], pp[620], r19c[11], r19s[12], r19c[12]);
FA	inst1596	(r18s[14], pp[590], r19c[12], r19s[13], r19c[13]);
FA	inst1597	(r18s[15], pp[591], r19c[13], r19s[14], r19c[14]);
FA	inst1598	(r18s[16], pp[592], r19c[14], r19s[15], r19c[15]);
FA	inst1599	(r18s[17], pp[593], r19c[15], r19s[16], r19c[16]);
FA	inst1600	(r18s[18], pp[594], r19c[16], r19s[17], r19c[17]);
FA	inst1601	(r18s[19], pp[595], r19c[17], r19s[18], r19c[18]);
FA	inst1602	(r18s[20], pp[596], r19c[18], r19s[19], r19c[19]);
FA	inst1603	(r18s[21], pp[597], r19c[19], r19s[20], r19c[20]);
FA	inst1604	(r18s[22], pp[598], r19c[20], r19s[21], r19c[21]);
FA	inst1605	(r18s[23], pp[599], r19c[21], r19s[22], r19c[22]);
FA	inst1606	(r18s[24], pp[600], r19c[22], r19s[23], r19c[23]);
FA	inst1607	(r18s[25], pp[601], r19c[23], r19s[24], r19c[24]);
FA	inst1608	(r18s[26], pp[602], r19c[24], r19s[25], r19c[25]);
FA	inst1609	(r18s[27], pp[603], r19c[25], r19s[26], r19c[26]);
FA	inst1610	(r18s[28], pp[604], r19c[26], r19s[27], r19c[27]);
FA	inst1611	(r18s[29], pp[605], r19c[27], r19s[28], r19c[28]);
FA	inst1612	(r18s[30], pp[606], r19c[28], r19s[29], r19c[29]);
FA	inst1613	(r18c[30], pp[607], r19c[29], r19s[30], r19c[30]);

HA	inst1614	(r19s[1], pp[640], m[20], r20c[0]);
FA	inst1615	(r19s[2], pp[641], r20c[0], r20s[1], r20c[1]);
FA	inst1616	(r19s[3], pp[642], r20c[1], r20s[2], r20c[2]);
FA	inst1617	(r19s[4], pp[643], r20c[2], r20s[3], r20c[3]);
FA	inst1618	(r19s[5], pp[644], r20c[3], r20s[4], r20c[4]);
FA	inst1619	(r19s[6], pp[645], r20c[4], r20s[5], r20c[5]);
FA	inst1620	(r19s[7], pp[646], r20c[5], r20s[6], r20c[6]);
FA	inst1621	(r19s[8], pp[647], r20c[6], r20s[7], r20c[7]);
FA	inst1622	(r19s[9], pp[648], r20c[7], r20s[8], r20c[8]);
FA	inst1623	(r19s[10], pp[649], r20c[8], r20s[9], r20c[9]);
FA	inst1624	(r19s[11], pp[650], r20c[9], r20s[10], r20c[10]);
FA	inst1625	(r19s[12], pp[651], r20c[10], r20s[11], r20c[11]);
FA	inst1626	(r19s[13], pp[621], r20c[11], r20s[12], r20c[12]);
FA	inst1627	(r19s[14], pp[622], r20c[12], r20s[13], r20c[13]);
FA	inst1628	(r19s[15], pp[623], r20c[13], r20s[14], r20c[14]);
FA	inst1629	(r19s[16], pp[624], r20c[14], r20s[15], r20c[15]);
FA	inst1630	(r19s[17], pp[625], r20c[15], r20s[16], r20c[16]);
FA	inst1631	(r19s[18], pp[626], r20c[16], r20s[17], r20c[17]);
FA	inst1632	(r19s[19], pp[627], r20c[17], r20s[18], r20c[18]);
FA	inst1633	(r19s[20], pp[628], r20c[18], r20s[19], r20c[19]);
FA	inst1634	(r19s[21], pp[629], r20c[19], r20s[20], r20c[20]);
FA	inst1635	(r19s[22], pp[630], r20c[20], r20s[21], r20c[21]);
FA	inst1636	(r19s[23], pp[631], r20c[21], r20s[22], r20c[22]);
FA	inst1637	(r19s[24], pp[632], r20c[22], r20s[23], r20c[23]);
FA	inst1638	(r19s[25], pp[633], r20c[23], r20s[24], r20c[24]);
FA	inst1639	(r19s[26], pp[634], r20c[24], r20s[25], r20c[25]);
FA	inst1640	(r19s[27], pp[635], r20c[25], r20s[26], r20c[26]);
FA	inst1641	(r19s[28], pp[636], r20c[26], r20s[27], r20c[27]);
FA	inst1642	(r19s[29], pp[637], r20c[27], r20s[28], r20c[28]);
FA	inst1643	(r19s[30], pp[638], r20c[28], r20s[29], r20c[29]);
FA	inst1644	(r19c[30], pp[639], r20c[29], r20s[30], r20c[30]);

HA	inst1645	(r20s[1], pp[672], m[21], r21c[0]);
FA	inst1646	(r20s[2], pp[673], r21c[0], r21s[1], r21c[1]);
FA	inst1647	(r20s[3], pp[674], r21c[1], r21s[2], r21c[2]);
FA	inst1648	(r20s[4], pp[675], r21c[2], r21s[3], r21c[3]);
FA	inst1649	(r20s[5], pp[676], r21c[3], r21s[4], r21c[4]);
FA	inst1650	(r20s[6], pp[677], r21c[4], r21s[5], r21c[5]);
FA	inst1651	(r20s[7], pp[678], r21c[5], r21s[6], r21c[6]);
FA	inst1652	(r20s[8], pp[679], r21c[6], r21s[7], r21c[7]);
FA	inst1653	(r20s[9], pp[680], r21c[7], r21s[8], r21c[8]);
FA	inst1654	(r20s[10], pp[681], r21c[8], r21s[9], r21c[9]);
FA	inst1655	(r20s[11], pp[682], r21c[9], r21s[10], r21c[10]);
FA	inst1656	(r20s[12], pp[652], r21c[10], r21s[11], r21c[11]);
FA	inst1657	(r20s[13], pp[653], r21c[11], r21s[12], r21c[12]);
FA	inst1658	(r20s[14], pp[654], r21c[12], r21s[13], r21c[13]);
FA	inst1659	(r20s[15], pp[655], r21c[13], r21s[14], r21c[14]);
FA	inst1660	(r20s[16], pp[656], r21c[14], r21s[15], r21c[15]);
FA	inst1661	(r20s[17], pp[657], r21c[15], r21s[16], r21c[16]);
FA	inst1662	(r20s[18], pp[658], r21c[16], r21s[17], r21c[17]);
FA	inst1663	(r20s[19], pp[659], r21c[17], r21s[18], r21c[18]);
FA	inst1664	(r20s[20], pp[660], r21c[18], r21s[19], r21c[19]);
FA	inst1665	(r20s[21], pp[661], r21c[19], r21s[20], r21c[20]);
FA	inst1666	(r20s[22], pp[662], r21c[20], r21s[21], r21c[21]);
FA	inst1667	(r20s[23], pp[663], r21c[21], r21s[22], r21c[22]);
FA	inst1668	(r20s[24], pp[664], r21c[22], r21s[23], r21c[23]);
FA	inst1669	(r20s[25], pp[665], r21c[23], r21s[24], r21c[24]);
FA	inst1670	(r20s[26], pp[666], r21c[24], r21s[25], r21c[25]);
FA	inst1671	(r20s[27], pp[667], r21c[25], r21s[26], r21c[26]);
FA	inst1672	(r20s[28], pp[668], r21c[26], r21s[27], r21c[27]);
FA	inst1673	(r20s[29], pp[669], r21c[27], r21s[28], r21c[28]);
FA	inst1674	(r20s[30], pp[670], r21c[28], r21s[29], r21c[29]);
FA	inst1675	(r20c[30], pp[671], r21c[29], r21s[30], r21c[30]);

HA	inst1676	(r21s[1], pp[704], m[22], r22c[0]);
FA	inst1677	(r21s[2], pp[705], r22c[0], r22s[1], r22c[1]);
FA	inst1678	(r21s[3], pp[706], r22c[1], r22s[2], r22c[2]);
FA	inst1679	(r21s[4], pp[707], r22c[2], r22s[3], r22c[3]);
FA	inst1680	(r21s[5], pp[708], r22c[3], r22s[4], r22c[4]);
FA	inst1681	(r21s[6], pp[709], r22c[4], r22s[5], r22c[5]);
FA	inst1682	(r21s[7], pp[710], r22c[5], r22s[6], r22c[6]);
FA	inst1683	(r21s[8], pp[711], r22c[6], r22s[7], r22c[7]);
FA	inst1684	(r21s[9], pp[712], r22c[7], r22s[8], r22c[8]);
FA	inst1685	(r21s[10], pp[713], r22c[8], r22s[9], r22c[9]);
FA	inst1686	(r21s[11], pp[683], r22c[9], r22s[10], r22c[10]);
FA	inst1687	(r21s[12], pp[684], r22c[10], r22s[11], r22c[11]);
FA	inst1688	(r21s[13], pp[685], r22c[11], r22s[12], r22c[12]);
FA	inst1689	(r21s[14], pp[686], r22c[12], r22s[13], r22c[13]);
FA	inst1690	(r21s[15], pp[687], r22c[13], r22s[14], r22c[14]);
FA	inst1691	(r21s[16], pp[688], r22c[14], r22s[15], r22c[15]);
FA	inst1692	(r21s[17], pp[689], r22c[15], r22s[16], r22c[16]);
FA	inst1693	(r21s[18], pp[690], r22c[16], r22s[17], r22c[17]);
FA	inst1694	(r21s[19], pp[691], r22c[17], r22s[18], r22c[18]);
FA	inst1695	(r21s[20], pp[692], r22c[18], r22s[19], r22c[19]);
FA	inst1696	(r21s[21], pp[693], r22c[19], r22s[20], r22c[20]);
FA	inst1697	(r21s[22], pp[694], r22c[20], r22s[21], r22c[21]);
FA	inst1698	(r21s[23], pp[695], r22c[21], r22s[22], r22c[22]);
FA	inst1699	(r21s[24], pp[696], r22c[22], r22s[23], r22c[23]);
FA	inst1700	(r21s[25], pp[697], r22c[23], r22s[24], r22c[24]);
FA	inst1701	(r21s[26], pp[698], r22c[24], r22s[25], r22c[25]);
FA	inst1702	(r21s[27], pp[699], r22c[25], r22s[26], r22c[26]);
FA	inst1703	(r21s[28], pp[700], r22c[26], r22s[27], r22c[27]);
FA	inst1704	(r21s[29], pp[701], r22c[27], r22s[28], r22c[28]);
FA	inst1705	(r21s[30], pp[702], r22c[28], r22s[29], r22c[29]);
FA	inst1706	(r21c[30], pp[703], r22c[29], r22s[30], r22c[30]);

HA	inst1707	(r22s[1], pp[736], m[23], r23c[0]);
FA	inst1708	(r22s[2], pp[737], r23c[0], r23s[1], r23c[1]);
FA	inst1709	(r22s[3], pp[738], r23c[1], r23s[2], r23c[2]);
FA	inst1710	(r22s[4], pp[739], r23c[2], r23s[3], r23c[3]);
FA	inst1711	(r22s[5], pp[740], r23c[3], r23s[4], r23c[4]);
FA	inst1712	(r22s[6], pp[741], r23c[4], r23s[5], r23c[5]);
FA	inst1713	(r22s[7], pp[742], r23c[5], r23s[6], r23c[6]);
FA	inst1714	(r22s[8], pp[743], r23c[6], r23s[7], r23c[7]);
FA	inst1715	(r22s[9], pp[744], r23c[7], r23s[8], r23c[8]);
FA	inst1716	(r22s[10], pp[714], r23c[8], r23s[9], r23c[9]);
FA	inst1717	(r22s[11], pp[715], r23c[9], r23s[10], r23c[10]);
FA	inst1718	(r22s[12], pp[716], r23c[10], r23s[11], r23c[11]);
FA	inst1719	(r22s[13], pp[717], r23c[11], r23s[12], r23c[12]);
FA	inst1720	(r22s[14], pp[718], r23c[12], r23s[13], r23c[13]);
FA	inst1721	(r22s[15], pp[719], r23c[13], r23s[14], r23c[14]);
FA	inst1722	(r22s[16], pp[720], r23c[14], r23s[15], r23c[15]);
FA	inst1723	(r22s[17], pp[721], r23c[15], r23s[16], r23c[16]);
FA	inst1724	(r22s[18], pp[722], r23c[16], r23s[17], r23c[17]);
FA	inst1725	(r22s[19], pp[723], r23c[17], r23s[18], r23c[18]);
FA	inst1726	(r22s[20], pp[724], r23c[18], r23s[19], r23c[19]);
FA	inst1727	(r22s[21], pp[725], r23c[19], r23s[20], r23c[20]);
FA	inst1728	(r22s[22], pp[726], r23c[20], r23s[21], r23c[21]);
FA	inst1729	(r22s[23], pp[727], r23c[21], r23s[22], r23c[22]);
FA	inst1730	(r22s[24], pp[728], r23c[22], r23s[23], r23c[23]);
FA	inst1731	(r22s[25], pp[729], r23c[23], r23s[24], r23c[24]);
FA	inst1732	(r22s[26], pp[730], r23c[24], r23s[25], r23c[25]);
FA	inst1733	(r22s[27], pp[731], r23c[25], r23s[26], r23c[26]);
FA	inst1734	(r22s[28], pp[732], r23c[26], r23s[27], r23c[27]);
FA	inst1735	(r22s[29], pp[733], r23c[27], r23s[28], r23c[28]);
FA	inst1736	(r22s[30], pp[734], r23c[28], r23s[29], r23c[29]);
FA	inst1737	(r22c[30], pp[735], r23c[29], r23s[30], r23c[30]);

HA	inst1738	(r23s[1], pp[768], m[24], r24c[0]);
FA	inst1739	(r23s[2], pp[769], r24c[0], r24s[1], r24c[1]);
FA	inst1740	(r23s[3], pp[770], r24c[1], r24s[2], r24c[2]);
FA	inst1741	(r23s[4], pp[771], r24c[2], r24s[3], r24c[3]);
FA	inst1742	(r23s[5], pp[772], r24c[3], r24s[4], r24c[4]);
FA	inst1743	(r23s[6], pp[773], r24c[4], r24s[5], r24c[5]);
FA	inst1744	(r23s[7], pp[774], r24c[5], r24s[6], r24c[6]);
FA	inst1745	(r23s[8], pp[775], r24c[6], r24s[7], r24c[7]);
FA	inst1746	(r23s[9], pp[745], r24c[7], r24s[8], r24c[8]);
FA	inst1747	(r23s[10], pp[746], r24c[8], r24s[9], r24c[9]);
FA	inst1748	(r23s[11], pp[747], r24c[9], r24s[10], r24c[10]);
FA	inst1749	(r23s[12], pp[748], r24c[10], r24s[11], r24c[11]);
FA	inst1750	(r23s[13], pp[749], r24c[11], r24s[12], r24c[12]);
FA	inst1751	(r23s[14], pp[750], r24c[12], r24s[13], r24c[13]);
FA	inst1752	(r23s[15], pp[751], r24c[13], r24s[14], r24c[14]);
FA	inst1753	(r23s[16], pp[752], r24c[14], r24s[15], r24c[15]);
FA	inst1754	(r23s[17], pp[753], r24c[15], r24s[16], r24c[16]);
FA	inst1755	(r23s[18], pp[754], r24c[16], r24s[17], r24c[17]);
FA	inst1756	(r23s[19], pp[755], r24c[17], r24s[18], r24c[18]);
FA	inst1757	(r23s[20], pp[756], r24c[18], r24s[19], r24c[19]);
FA	inst1758	(r23s[21], pp[757], r24c[19], r24s[20], r24c[20]);
FA	inst1759	(r23s[22], pp[758], r24c[20], r24s[21], r24c[21]);
FA	inst1760	(r23s[23], pp[759], r24c[21], r24s[22], r24c[22]);
FA	inst1761	(r23s[24], pp[760], r24c[22], r24s[23], r24c[23]);
FA	inst1762	(r23s[25], pp[761], r24c[23], r24s[24], r24c[24]);
FA	inst1763	(r23s[26], pp[762], r24c[24], r24s[25], r24c[25]);
FA	inst1764	(r23s[27], pp[763], r24c[25], r24s[26], r24c[26]);
FA	inst1765	(r23s[28], pp[764], r24c[26], r24s[27], r24c[27]);
FA	inst1766	(r23s[29], pp[765], r24c[27], r24s[28], r24c[28]);
FA	inst1767	(r23s[30], pp[766], r24c[28], r24s[29], r24c[29]);
FA	inst1768	(r23c[30], pp[767], r24c[29], r24s[30], r24c[30]);

HA	inst1769	(r24s[1], pp[800], m[25], r25c[0]);
FA	inst1770	(r24s[2], pp[801], r25c[0], r25s[1], r25c[1]);
FA	inst1771	(r24s[3], pp[802], r25c[1], r25s[2], r25c[2]);
FA	inst1772	(r24s[4], pp[803], r25c[2], r25s[3], r25c[3]);
FA	inst1773	(r24s[5], pp[804], r25c[3], r25s[4], r25c[4]);
FA	inst1774	(r24s[6], pp[805], r25c[4], r25s[5], r25c[5]);
FA	inst1775	(r24s[7], pp[806], r25c[5], r25s[6], r25c[6]);
FA	inst1776	(r24s[8], pp[776], r25c[6], r25s[7], r25c[7]);
FA	inst1777	(r24s[9], pp[777], r25c[7], r25s[8], r25c[8]);
FA	inst1778	(r24s[10], pp[778], r25c[8], r25s[9], r25c[9]);
FA	inst1779	(r24s[11], pp[779], r25c[9], r25s[10], r25c[10]);
FA	inst1780	(r24s[12], pp[780], r25c[10], r25s[11], r25c[11]);
FA	inst1781	(r24s[13], pp[781], r25c[11], r25s[12], r25c[12]);
FA	inst1782	(r24s[14], pp[782], r25c[12], r25s[13], r25c[13]);
FA	inst1783	(r24s[15], pp[783], r25c[13], r25s[14], r25c[14]);
FA	inst1784	(r24s[16], pp[784], r25c[14], r25s[15], r25c[15]);
FA	inst1785	(r24s[17], pp[785], r25c[15], r25s[16], r25c[16]);
FA	inst1786	(r24s[18], pp[786], r25c[16], r25s[17], r25c[17]);
FA	inst1787	(r24s[19], pp[787], r25c[17], r25s[18], r25c[18]);
FA	inst1788	(r24s[20], pp[788], r25c[18], r25s[19], r25c[19]);
FA	inst1789	(r24s[21], pp[789], r25c[19], r25s[20], r25c[20]);
FA	inst1790	(r24s[22], pp[790], r25c[20], r25s[21], r25c[21]);
FA	inst1791	(r24s[23], pp[791], r25c[21], r25s[22], r25c[22]);
FA	inst1792	(r24s[24], pp[792], r25c[22], r25s[23], r25c[23]);
FA	inst1793	(r24s[25], pp[793], r25c[23], r25s[24], r25c[24]);
FA	inst1794	(r24s[26], pp[794], r25c[24], r25s[25], r25c[25]);
FA	inst1795	(r24s[27], pp[795], r25c[25], r25s[26], r25c[26]);
FA	inst1796	(r24s[28], pp[796], r25c[26], r25s[27], r25c[27]);
FA	inst1797	(r24s[29], pp[797], r25c[27], r25s[28], r25c[28]);
FA	inst1798	(r24s[30], pp[798], r25c[28], r25s[29], r25c[29]);
FA	inst1799	(r24c[30], pp[799], r25c[29], r25s[30], r25c[30]);

HA	inst1800	(r25s[1], pp[832], m[26], r26c[0]);
FA	inst1801	(r25s[2], pp[833], r26c[0], r26s[1], r26c[1]);
FA	inst1802	(r25s[3], pp[834], r26c[1], r26s[2], r26c[2]);
FA	inst1803	(r25s[4], pp[835], r26c[2], r26s[3], r26c[3]);
FA	inst1804	(r25s[5], pp[836], r26c[3], r26s[4], r26c[4]);
FA	inst1805	(r25s[6], pp[837], r26c[4], r26s[5], r26c[5]);
FA	inst1806	(r25s[7], pp[807], r26c[5], r26s[6], r26c[6]);
FA	inst1807	(r25s[8], pp[808], r26c[6], r26s[7], r26c[7]);
FA	inst1808	(r25s[9], pp[809], r26c[7], r26s[8], r26c[8]);
FA	inst1809	(r25s[10], pp[810], r26c[8], r26s[9], r26c[9]);
FA	inst1810	(r25s[11], pp[811], r26c[9], r26s[10], r26c[10]);
FA	inst1811	(r25s[12], pp[812], r26c[10], r26s[11], r26c[11]);
FA	inst1812	(r25s[13], pp[813], r26c[11], r26s[12], r26c[12]);
FA	inst1813	(r25s[14], pp[814], r26c[12], r26s[13], r26c[13]);
FA	inst1814	(r25s[15], pp[815], r26c[13], r26s[14], r26c[14]);
FA	inst1815	(r25s[16], pp[816], r26c[14], r26s[15], r26c[15]);
FA	inst1816	(r25s[17], pp[817], r26c[15], r26s[16], r26c[16]);
FA	inst1817	(r25s[18], pp[818], r26c[16], r26s[17], r26c[17]);
FA	inst1818	(r25s[19], pp[819], r26c[17], r26s[18], r26c[18]);
FA	inst1819	(r25s[20], pp[820], r26c[18], r26s[19], r26c[19]);
FA	inst1820	(r25s[21], pp[821], r26c[19], r26s[20], r26c[20]);
FA	inst1821	(r25s[22], pp[822], r26c[20], r26s[21], r26c[21]);
FA	inst1822	(r25s[23], pp[823], r26c[21], r26s[22], r26c[22]);
FA	inst1823	(r25s[24], pp[824], r26c[22], r26s[23], r26c[23]);
FA	inst1824	(r25s[25], pp[825], r26c[23], r26s[24], r26c[24]);
FA	inst1825	(r25s[26], pp[826], r26c[24], r26s[25], r26c[25]);
FA	inst1826	(r25s[27], pp[827], r26c[25], r26s[26], r26c[26]);
FA	inst1827	(r25s[28], pp[828], r26c[26], r26s[27], r26c[27]);
FA	inst1828	(r25s[29], pp[829], r26c[27], r26s[28], r26c[28]);
FA	inst1829	(r25s[30], pp[830], r26c[28], r26s[29], r26c[29]);
FA	inst1830	(r25c[30], pp[831], r26c[29], r26s[30], r26c[30]);

HA	inst1831	(r26s[1], pp[864], m[27], r27c[0]);
FA	inst1832	(r26s[2], pp[865], r27c[0], r27s[1], r27c[1]);
FA	inst1833	(r26s[3], pp[866], r27c[1], r27s[2], r27c[2]);
FA	inst1834	(r26s[4], pp[867], r27c[2], r27s[3], r27c[3]);
FA	inst1835	(r26s[5], pp[868], r27c[3], r27s[4], r27c[4]);
FA	inst1836	(r26s[6], pp[838], r27c[4], r27s[5], r27c[5]);
FA	inst1837	(r26s[7], pp[839], r27c[5], r27s[6], r27c[6]);
FA	inst1838	(r26s[8], pp[840], r27c[6], r27s[7], r27c[7]);
FA	inst1839	(r26s[9], pp[841], r27c[7], r27s[8], r27c[8]);
FA	inst1840	(r26s[10], pp[842], r27c[8], r27s[9], r27c[9]);
FA	inst1841	(r26s[11], pp[843], r27c[9], r27s[10], r27c[10]);
FA	inst1842	(r26s[12], pp[844], r27c[10], r27s[11], r27c[11]);
FA	inst1843	(r26s[13], pp[845], r27c[11], r27s[12], r27c[12]);
FA	inst1844	(r26s[14], pp[846], r27c[12], r27s[13], r27c[13]);
FA	inst1845	(r26s[15], pp[847], r27c[13], r27s[14], r27c[14]);
FA	inst1846	(r26s[16], pp[848], r27c[14], r27s[15], r27c[15]);
FA	inst1847	(r26s[17], pp[849], r27c[15], r27s[16], r27c[16]);
FA	inst1848	(r26s[18], pp[850], r27c[16], r27s[17], r27c[17]);
FA	inst1849	(r26s[19], pp[851], r27c[17], r27s[18], r27c[18]);
FA	inst1850	(r26s[20], pp[852], r27c[18], r27s[19], r27c[19]);
FA	inst1851	(r26s[21], pp[853], r27c[19], r27s[20], r27c[20]);
FA	inst1852	(r26s[22], pp[854], r27c[20], r27s[21], r27c[21]);
FA	inst1853	(r26s[23], pp[855], r27c[21], r27s[22], r27c[22]);
FA	inst1854	(r26s[24], pp[856], r27c[22], r27s[23], r27c[23]);
FA	inst1855	(r26s[25], pp[857], r27c[23], r27s[24], r27c[24]);
FA	inst1856	(r26s[26], pp[858], r27c[24], r27s[25], r27c[25]);
FA	inst1857	(r26s[27], pp[859], r27c[25], r27s[26], r27c[26]);
FA	inst1858	(r26s[28], pp[860], r27c[26], r27s[27], r27c[27]);
FA	inst1859	(r26s[29], pp[861], r27c[27], r27s[28], r27c[28]);
FA	inst1860	(r26s[30], pp[862], r27c[28], r27s[29], r27c[29]);
FA	inst1861	(r26c[30], pp[863], r27c[29], r27s[30], r27c[30]);

HA	inst1862	(r27s[1], pp[896], m[28], r28c[0]);
FA	inst1863	(r27s[2], pp[897], r28c[0], r28s[1], r28c[1]);
FA	inst1864	(r27s[3], pp[898], r28c[1], r28s[2], r28c[2]);
FA	inst1865	(r27s[4], pp[899], r28c[2], r28s[3], r28c[3]);
FA	inst1866	(r27s[5], pp[869], r28c[3], r28s[4], r28c[4]);
FA	inst1867	(r27s[6], pp[870], r28c[4], r28s[5], r28c[5]);
FA	inst1868	(r27s[7], pp[871], r28c[5], r28s[6], r28c[6]);
FA	inst1869	(r27s[8], pp[872], r28c[6], r28s[7], r28c[7]);
FA	inst1870	(r27s[9], pp[873], r28c[7], r28s[8], r28c[8]);
FA	inst1871	(r27s[10], pp[874], r28c[8], r28s[9], r28c[9]);
FA	inst1872	(r27s[11], pp[875], r28c[9], r28s[10], r28c[10]);
FA	inst1873	(r27s[12], pp[876], r28c[10], r28s[11], r28c[11]);
FA	inst1874	(r27s[13], pp[877], r28c[11], r28s[12], r28c[12]);
FA	inst1875	(r27s[14], pp[878], r28c[12], r28s[13], r28c[13]);
FA	inst1876	(r27s[15], pp[879], r28c[13], r28s[14], r28c[14]);
FA	inst1877	(r27s[16], pp[880], r28c[14], r28s[15], r28c[15]);
FA	inst1878	(r27s[17], pp[881], r28c[15], r28s[16], r28c[16]);
FA	inst1879	(r27s[18], pp[882], r28c[16], r28s[17], r28c[17]);
FA	inst1880	(r27s[19], pp[883], r28c[17], r28s[18], r28c[18]);
FA	inst1881	(r27s[20], pp[884], r28c[18], r28s[19], r28c[19]);
FA	inst1882	(r27s[21], pp[885], r28c[19], r28s[20], r28c[20]);
FA	inst1883	(r27s[22], pp[886], r28c[20], r28s[21], r28c[21]);
FA	inst1884	(r27s[23], pp[887], r28c[21], r28s[22], r28c[22]);
FA	inst1885	(r27s[24], pp[888], r28c[22], r28s[23], r28c[23]);
FA	inst1886	(r27s[25], pp[889], r28c[23], r28s[24], r28c[24]);
FA	inst1887	(r27s[26], pp[890], r28c[24], r28s[25], r28c[25]);
FA	inst1888	(r27s[27], pp[891], r28c[25], r28s[26], r28c[26]);
FA	inst1889	(r27s[28], pp[892], r28c[26], r28s[27], r28c[27]);
FA	inst1890	(r27s[29], pp[893], r28c[27], r28s[28], r28c[28]);
FA	inst1891	(r27s[30], pp[894], r28c[28], r28s[29], r28c[29]);
FA	inst1892	(r27c[30], pp[895], r28c[29], r28s[30], r28c[30]);

HA	inst1893	(r28s[1], pp[928], m[29], r29c[0]);
FA	inst1894	(r28s[2], pp[929], r29c[0], r29s[1], r29c[1]);
FA	inst1895	(r28s[3], pp[930], r29c[1], r29s[2], r29c[2]);
FA	inst1896	(r28s[4], pp[900], r29c[2], r29s[3], r29c[3]);
FA	inst1897	(r28s[5], pp[901], r29c[3], r29s[4], r29c[4]);
FA	inst1898	(r28s[6], pp[902], r29c[4], r29s[5], r29c[5]);
FA	inst1899	(r28s[7], pp[903], r29c[5], r29s[6], r29c[6]);
FA	inst1900	(r28s[8], pp[904], r29c[6], r29s[7], r29c[7]);
FA	inst1901	(r28s[9], pp[905], r29c[7], r29s[8], r29c[8]);
FA	inst1902	(r28s[10], pp[906], r29c[8], r29s[9], r29c[9]);
FA	inst1903	(r28s[11], pp[907], r29c[9], r29s[10], r29c[10]);
FA	inst1904	(r28s[12], pp[908], r29c[10], r29s[11], r29c[11]);
FA	inst1905	(r28s[13], pp[909], r29c[11], r29s[12], r29c[12]);
FA	inst1906	(r28s[14], pp[910], r29c[12], r29s[13], r29c[13]);
FA	inst1907	(r28s[15], pp[911], r29c[13], r29s[14], r29c[14]);
FA	inst1908	(r28s[16], pp[912], r29c[14], r29s[15], r29c[15]);
FA	inst1909	(r28s[17], pp[913], r29c[15], r29s[16], r29c[16]);
FA	inst1910	(r28s[18], pp[914], r29c[16], r29s[17], r29c[17]);
FA	inst1911	(r28s[19], pp[915], r29c[17], r29s[18], r29c[18]);
FA	inst1912	(r28s[20], pp[916], r29c[18], r29s[19], r29c[19]);
FA	inst1913	(r28s[21], pp[917], r29c[19], r29s[20], r29c[20]);
FA	inst1914	(r28s[22], pp[918], r29c[20], r29s[21], r29c[21]);
FA	inst1915	(r28s[23], pp[919], r29c[21], r29s[22], r29c[22]);
FA	inst1916	(r28s[24], pp[920], r29c[22], r29s[23], r29c[23]);
FA	inst1917	(r28s[25], pp[921], r29c[23], r29s[24], r29c[24]);
FA	inst1918	(r28s[26], pp[922], r29c[24], r29s[25], r29c[25]);
FA	inst1919	(r28s[27], pp[923], r29c[25], r29s[26], r29c[26]);
FA	inst1920	(r28s[28], pp[924], r29c[26], r29s[27], r29c[27]);
FA	inst1921	(r28s[29], pp[925], r29c[27], r29s[28], r29c[28]);
FA	inst1922	(r28s[30], pp[926], r29c[28], r29s[29], r29c[29]);
FA	inst1923	(r28c[30], pp[927], r29c[29], r29s[30], r29c[30]);

HA	inst1924	(r29s[1], pp[960], m[30], r30c[0]);
FA	inst1925	(r29s[2], pp[961], r30c[0], r30s[1], r30c[1]);
FA	inst1926	(r29s[3], pp[931], r30c[1], r30s[2], r30c[2]);
FA	inst1927	(r29s[4], pp[932], r30c[2], r30s[3], r30c[3]);
FA	inst1928	(r29s[5], pp[933], r30c[3], r30s[4], r30c[4]);
FA	inst1929	(r29s[6], pp[934], r30c[4], r30s[5], r30c[5]);
FA	inst1930	(r29s[7], pp[935], r30c[5], r30s[6], r30c[6]);
FA	inst1931	(r29s[8], pp[936], r30c[6], r30s[7], r30c[7]);
FA	inst1932	(r29s[9], pp[937], r30c[7], r30s[8], r30c[8]);
FA	inst1933	(r29s[10], pp[938], r30c[8], r30s[9], r30c[9]);
FA	inst1934	(r29s[11], pp[939], r30c[9], r30s[10], r30c[10]);
FA	inst1935	(r29s[12], pp[940], r30c[10], r30s[11], r30c[11]);
FA	inst1936	(r29s[13], pp[941], r30c[11], r30s[12], r30c[12]);
FA	inst1937	(r29s[14], pp[942], r30c[12], r30s[13], r30c[13]);
FA	inst1938	(r29s[15], pp[943], r30c[13], r30s[14], r30c[14]);
FA	inst1939	(r29s[16], pp[944], r30c[14], r30s[15], r30c[15]);
FA	inst1940	(r29s[17], pp[945], r30c[15], r30s[16], r30c[16]);
FA	inst1941	(r29s[18], pp[946], r30c[16], r30s[17], r30c[17]);
FA	inst1942	(r29s[19], pp[947], r30c[17], r30s[18], r30c[18]);
FA	inst1943	(r29s[20], pp[948], r30c[18], r30s[19], r30c[19]);
FA	inst1944	(r29s[21], pp[949], r30c[19], r30s[20], r30c[20]);
FA	inst1945	(r29s[22], pp[950], r30c[20], r30s[21], r30c[21]);
FA	inst1946	(r29s[23], pp[951], r30c[21], r30s[22], r30c[22]);
FA	inst1947	(r29s[24], pp[952], r30c[22], r30s[23], r30c[23]);
FA	inst1948	(r29s[25], pp[953], r30c[23], r30s[24], r30c[24]);
FA	inst1949	(r29s[26], pp[954], r30c[24], r30s[25], r30c[25]);
FA	inst1950	(r29s[27], pp[955], r30c[25], r30s[26], r30c[26]);
FA	inst1951	(r29s[28], pp[956], r30c[26], r30s[27], r30c[27]);
FA	inst1952	(r29s[29], pp[957], r30c[27], r30s[28], r30c[28]);
FA	inst1953	(r29s[30], pp[958], r30c[28], r30s[29], r30c[29]);
FA	inst1954	(r29c[30], pp[959], r30c[29], r30s[30], r30c[30]);

HA	inst1955	(r30s[1], pp[992], m[31], r31c[0]);
FA	inst1956	(r30s[2], pp[962], r31c[0], r31s[1], r31c[1]);
FA	inst1957	(r30s[3], pp[963], r31c[1], r31s[2], r31c[2]);
FA	inst1958	(r30s[4], pp[964], r31c[2], r31s[3], r31c[3]);
FA	inst1959	(r30s[5], pp[965], r31c[3], r31s[4], r31c[4]);
FA	inst1960	(r30s[6], pp[966], r31c[4], r31s[5], r31c[5]);
FA	inst1961	(r30s[7], pp[967], r31c[5], r31s[6], r31c[6]);
FA	inst1962	(r30s[8], pp[968], r31c[6], r31s[7], r31c[7]);
FA	inst1963	(r30s[9], pp[969], r31c[7], r31s[8], r31c[8]);
FA	inst1964	(r30s[10], pp[970], r31c[8], r31s[9], r31c[9]);
FA	inst1965	(r30s[11], pp[971], r31c[9], r31s[10], r31c[10]);
FA	inst1966	(r30s[12], pp[972], r31c[10], r31s[11], r31c[11]);
FA	inst1967	(r30s[13], pp[973], r31c[11], r31s[12], r31c[12]);
FA	inst1968	(r30s[14], pp[974], r31c[12], r31s[13], r31c[13]);
FA	inst1969	(r30s[15], pp[975], r31c[13], r31s[14], r31c[14]);
FA	inst1970	(r30s[16], pp[976], r31c[14], r31s[15], r31c[15]);
FA	inst1971	(r30s[17], pp[977], r31c[15], r31s[16], r31c[16]);
FA	inst1972	(r30s[18], pp[978], r31c[16], r31s[17], r31c[17]);
FA	inst1973	(r30s[19], pp[979], r31c[17], r31s[18], r31c[18]);
FA	inst1974	(r30s[20], pp[980], r31c[18], r31s[19], r31c[19]);
FA	inst1975	(r30s[21], pp[981], r31c[19], r31s[20], r31c[20]);
FA	inst1976	(r30s[22], pp[982], r31c[20], r31s[21], r31c[21]);
FA	inst1977	(r30s[23], pp[983], r31c[21], r31s[22], r31c[22]);
FA	inst1978	(r30s[24], pp[984], r31c[22], r31s[23], r31c[23]);
FA	inst1979	(r30s[25], pp[985], r31c[23], r31s[24], r31c[24]);
FA	inst1980	(r30s[26], pp[986], r31c[24], r31s[25], r31c[25]);
FA	inst1981	(r30s[27], pp[987], r31c[25], r31s[26], r31c[26]);
FA	inst1982	(r30s[28], pp[988], r31c[26], r31s[27], r31c[27]);
FA	inst1983	(r30s[29], pp[989], r31c[27], r31s[28], r31c[28]);
FA	inst1984	(r30s[30], pp[990], r31c[28], r31s[29], r31c[29]);
FA	inst1985	(r30c[30], pp[991], r31c[29], r31s[30], r31c[30]);

HA	inst1986	(r31s[1], pp[993], m[32], r32c[0]);
FA	inst1987	(r31s[2], pp[994], r32c[0], m[33], r32c[1]);
FA	inst1988	(r31s[3], pp[995], r32c[1], m[34], r32c[2]);
FA	inst1989	(r31s[4], pp[996], r32c[2], m[35], r32c[3]);
FA	inst1990	(r31s[5], pp[997], r32c[3], m[36], r32c[4]);
FA	inst1991	(r31s[6], pp[998], r32c[4], m[37], r32c[5]);
FA	inst1992	(r31s[7], pp[999], r32c[5], m[38], r32c[6]);
FA	inst1993	(r31s[8], pp[1000], r32c[6], m[39], r32c[7]);
FA	inst1994	(r31s[9], pp[1001], r32c[7], m[40], r32c[8]);
FA	inst1995	(r31s[10], pp[1002], r32c[8], m[41], r32c[9]);
FA	inst1996	(r31s[11], pp[1003], r32c[9], m[42], r32c[10]);
FA	inst1997	(r31s[12], pp[1004], r32c[10], m[43], r32c[11]);
FA	inst1998	(r31s[13], pp[1005], r32c[11], m[44], r32c[12]);
FA	inst1999	(r31s[14], pp[1006], r32c[12], m[45], r32c[13]);
FA	inst2000	(r31s[15], pp[1007], r32c[13], m[46], r32c[14]);
FA	inst2001	(r31s[16], pp[1008], r32c[14], m[47], r32c[15]);
FA	inst2002	(r31s[17], pp[1009], r32c[15], m[48], r32c[16]);
FA	inst2003	(r31s[18], pp[1010], r32c[16], m[49], r32c[17]);
FA	inst2004	(r31s[19], pp[1011], r32c[17], m[50], r32c[18]);
FA	inst2005	(r31s[20], pp[1012], r32c[18], m[51], r32c[19]);
FA	inst2006	(r31s[21], pp[1013], r32c[19], m[52], r32c[20]);
FA	inst2007	(r31s[22], pp[1014], r32c[20], m[53], r32c[21]);
FA	inst2008	(r31s[23], pp[1015], r32c[21], m[54], r32c[22]);
FA	inst2009	(r31s[24], pp[1016], r32c[22], m[55], r32c[23]);
FA	inst2010	(r31s[25], pp[1017], r32c[23], m[56], r32c[24]);
FA	inst2011	(r31s[26], pp[1018], r32c[24], m[57], r32c[25]);
FA	inst2012	(r31s[27], pp[1019], r32c[25], m[58], r32c[26]);
FA	inst2013	(r31s[28], pp[1020], r32c[26], m[59], r32c[27]);
FA	inst2014	(r31s[29], pp[1021], r32c[27], m[60], r32c[28]);
FA	inst2015	(r31s[30], pp[1022], r32c[28], m[61], r32c[29]);
FA	inst2016	(r31c[30], pp[1023], r32c[29], m[62], m[63]);
endmodule
