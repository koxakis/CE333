////////////////////////////////////////////////////////////////////////////////////
//Module name: Memory Controller Module
//File name: mem_ctrl.h
//Descreption: Provides control signals for memory modules 
////////////////////////////////////////////////////////////////////////////////////
module mem_ctrl(
	mc_clk,
	mc_reset,
	mc_data_address_in,
	mc_address_mem,
	mc_data_in,
	mc_data_out,
	mem_data_in,
	mem_data_out, 
	mc_data_contition,
	mc_err
);

endmodule // 