`timescale 1ns/10ps
module alu(
    clk,
	reset,
    inA,
    inB,
    opcode,
    result,
    extra_result,
    //zero,
    PStart,
    PDone
    );
    
    parameter ADD = 3'b000; //0
    parameter SUB = 3'b001; //1
    parameter OR  = 3'b010; //2
    parameter AND = 3'b011; //3
    parameter NOT = 3'b100; //4
    parameter MUL = 3'b101; //5
    parameter SLL = 3'b110; //6
    parameter SLR = 3'b111; //7
    
    input	clk, reset;
    input       [31:0]         inA, inB;
    input       [2:0]          opcode;
    output reg  [31:0]         result, extra_result;
    input wire                 PStart;
    output reg                 PDone; 
    
    reg [63:0]     total_result;
    wire[63:0]     mul_res;
    
    reg [31:0] inA_Reg, inB_Reg;
    reg [2:0] opcode_reg;
    reg ProcConditon_reg, ProcConditon_reg2;
	wire Pdone_out;

	wire o1, o2, xout;
    
    multiplier mu0(clk, inA_Reg, inB_Reg, mul_res, ProcConditon_reg, Pdone_out);

    
    always@(posedge clk or posedge reset)
    begin
	if (reset) begin
		PDone <= 1'b0;
		total_result = 64'b0;
		result <= 'b0;
		extra_result <= 'b0;
		ProcConditon_reg <='b0;

		inA_Reg <= 'b0;
		inB_Reg <= 'b0;
		opcode_reg <= 'b0;

	end else begin

		if (PStart) begin
	    	inA_Reg <= inA;
        	inB_Reg <= inB;
        	ProcConditon_reg <= PStart;
        	opcode_reg <= opcode;
			if (opcode_reg == MUL) begin
				PDone <= Pdone_out;
			end else begin
				PDone <= ProcConditon_reg;
			end
		end else begin
			ProcConditon_reg <= 1'b0;
		end
		    
        total_result = 64'b0;
    
        case(opcode_reg)
                ADD:
                begin
                    total_result = inA_Reg + inB_Reg;
                end
                
                SUB:
                begin
                    total_result = inA_Reg - inB_Reg;
                end
                
                OR:
                begin
                    total_result = inA_Reg | inB_Reg;
                end
                
                AND:
                begin
                    total_result = inA_Reg & inB_Reg;
                end
                
                NOT:
                begin
                    total_result = ~ inA_Reg;
                end
                
                MUL:
                begin
                    total_result = mul_res;
                end
                
                SLL:
                begin
                    total_result = inA_Reg << inB_Reg[4:0];
                end 
                
                SLR:
                begin
                    total_result = inA_Reg >> inB_Reg[4:0];
                end 
        endcase
        
        	result       <= total_result[ 31:0];
        	extra_result <= total_result[63:32];

		end 
	end
endmodule

module HA (I1, I2, sum, carry);
input I1, I2;
output sum, carry;
xor (sum, I1, I2);
and (carry, I1, I2);
endmodule

module FA (I1, I2, I3, sum, carry);
input I1, I2, I3;
output sum, carry;
wire o1, o2, xout;
xor (xout, I1, I2);
xor (sum, xout, I3);
and (o1, I1, I2);
and (o2, xout, I3);
or (carry, o1, o2);
endmodule

module multiplier (clk, a, b, m, PDone_in, PDone_out);
input clk;
input PDone_in;
output reg PDone_out;
input	[31 :0] a;
input	[31 :0] b;
output	[63 :0] m;

reg [31:0] ProcConditon_reg;

//reg ProcConditon_reg, ProcConditon_reg2, ProcConditon_reg3, ProcConditon_reg4, ProcConditon_reg5;
//reg ProcConditon_reg6, ProcConditon_reg7;


wire	[1023 :1]	pp;
reg     [1023 :1]   pp_reg; 
wire	[30 :0]	r1c;
wire	[30 :1]	r1s;
reg		[30 :1] r1s_reg;
reg		[30 :1] r23s_reg;
reg		[30 :1] r10s_reg;
reg		[31:0]  rc_last_reg;
wire	[30 :0]	r2c;
wire	[30 :1]	r2s;
reg		[30 :1] r2s_reg;
wire	[30 :0]	r3c;
wire	[30 :1]	r3s;
reg		[30 :1] r3s_reg;
wire	[30 :0]	r4c;
wire	[30 :1]	r4s;
reg		[30 :1] r4s_reg;
wire	[30 :0]	r5c;
reg		[30 :1] r5s_reg;
wire	[30 :1]	r5s;
wire	[30 :0]	r6c;
reg		[30 :1] r6s_reg;
wire	[30 :1]	r6s;
wire	[30 :0]	r7c;
reg		[30 :1] r7s_reg;
wire	[30 :1]	r7s;
wire	[30 :0]	r8c;
reg		[30 :1] r8s_reg;
wire	[30 :1]	r8s;
wire	[30 :0]	r9c;
reg		[30 :1] r9s_reg;
wire	[30 :1]	r9s;
wire	[30 :0]	r10c;
wire	[30 :1]	r10s;
wire	[30 :0]	r11c;
reg		[30 :1] r11s_reg;
wire	[30 :1]	r11s;
wire	[30 :0]	r12c;
reg		[30 :1] r12s_reg;
wire	[30 :1]	r12s;
wire	[30 :0]	r13c;
reg		[30 :1] r13s_reg;
wire	[30 :1]	r13s;
wire	[30 :0]	r14c;
reg		[30 :1] r14s_reg;
wire	[30 :1]	r14s;
wire	[30 :0]	r15c;
reg		[30 :1] r15s_reg;
wire	[30 :1]	r15s;
wire	[30 :0]	r16c;
reg		[30 :1] r16s_reg;
wire	[30 :1]	r16s;
wire	[30 :0]	r17c;
reg		[30 :1] r17s_reg;
wire	[30 :1]	r17s;
reg		[30 :1] r18s_reg;
wire	[30 :0]	r18c;
wire	[30 :1]	r18s;
reg		[30 :1] r19s_reg;
wire	[30 :0]	r19c;
wire	[30 :1]	r19s;
reg		[30 :1] r20s_reg;
wire	[30 :0]	r20c;
wire	[30 :1]	r20s;
reg		[30 :1] r21s_reg;
wire	[30 :0]	r21c;
wire	[30 :1]	r21s;
reg		[30 :1] r22s_reg;
wire	[30 :0]	r22c;
wire	[30 :1]	r22s;
wire	[30 :0]	r23c;
wire	[30 :1]	r23s;
reg		[30 :1] r24s_reg;
wire	[30 :0]	r24c;
wire	[30 :1]	r24s;
reg		[30 :1] r25s_reg;
wire	[30 :0]	r25c;
wire	[30 :1]	r25s;
reg		[30 :1] r26s_reg;
wire	[30 :0]	r26c;
wire	[30 :1]	r26s;
reg		[30 :1] r27s_reg;
wire	[30 :0]	r27c;
wire	[30 :1]	r27s;
reg		[30 :1] r28s_reg;
wire	[30 :0]	r28c;
wire	[30 :1]	r28s;
wire	[30 :0]	r29c;
reg		[30 :1] r29s_reg;
wire	[30 :1]	r29s;
wire	[30 :0]	r30c;
reg		[30 :1] r30s_reg;
wire	[30 :1]	r30s;
wire	[30 :0]	r31c;
reg		[30 :1] r31s_reg;
wire	[30 :1]	r31s;
wire	[29 :0]	r32c;

and	(m[0], a[0], b[0]);
and	(pp[1], a[0], b[1]);
and	(pp[2], a[0], b[2]);
and	(pp[3], a[0], b[3]);
and	(pp[4], a[0], b[4]);
and	(pp[5], a[0], b[5]);
and	(pp[6], a[0], b[6]);
and	(pp[7], a[0], b[7]);
and	(pp[8], a[0], b[8]);
and	(pp[9], a[0], b[9]);
and	(pp[10], a[0], b[10]);
and	(pp[11], a[0], b[11]);
and	(pp[12], a[0], b[12]);
and	(pp[13], a[0], b[13]);
and	(pp[14], a[0], b[14]);
and	(pp[15], a[0], b[15]);
and	(pp[16], a[0], b[16]);
and	(pp[17], a[0], b[17]);
and	(pp[18], a[0], b[18]);
and	(pp[19], a[0], b[19]);
and	(pp[20], a[0], b[20]);
and	(pp[21], a[0], b[21]);
and	(pp[22], a[0], b[22]);
and	(pp[23], a[0], b[23]);
and	(pp[24], a[0], b[24]);
and	(pp[25], a[0], b[25]);
and	(pp[26], a[0], b[26]);
and	(pp[27], a[0], b[27]);
and	(pp[28], a[0], b[28]);
and	(pp[29], a[0], b[29]);
and	(pp[30], a[0], b[30]);
and	(pp[31], a[0], b[31]);
and	(pp[32], a[1], b[0]);
and	(pp[33], a[1], b[1]);
and	(pp[34], a[1], b[2]);
and	(pp[35], a[1], b[3]);
and	(pp[36], a[1], b[4]);
and	(pp[37], a[1], b[5]);
and	(pp[38], a[1], b[6]);
and	(pp[39], a[1], b[7]);
and	(pp[40], a[1], b[8]);
and	(pp[41], a[1], b[9]);
and	(pp[42], a[1], b[10]);
and	(pp[43], a[1], b[11]);
and	(pp[44], a[1], b[12]);
and	(pp[45], a[1], b[13]);
and	(pp[46], a[1], b[14]);
and	(pp[47], a[1], b[15]);
and	(pp[48], a[1], b[16]);
and	(pp[49], a[1], b[17]);
and	(pp[50], a[1], b[18]);
and	(pp[51], a[1], b[19]);
and	(pp[52], a[1], b[20]);
and	(pp[53], a[1], b[21]);
and	(pp[54], a[1], b[22]);
and	(pp[55], a[1], b[23]);
and	(pp[56], a[1], b[24]);
and	(pp[57], a[1], b[25]);
and	(pp[58], a[1], b[26]);
and	(pp[59], a[1], b[27]);
and	(pp[60], a[1], b[28]);
and	(pp[61], a[1], b[29]);
and	(pp[62], a[1], b[30]);
and	(pp[63], a[1], b[31]);
and	(pp[64], a[2], b[0]);
and	(pp[65], a[2], b[1]);
and	(pp[66], a[2], b[2]);
and	(pp[67], a[2], b[3]);
and	(pp[68], a[2], b[4]);
and	(pp[69], a[2], b[5]);
and	(pp[70], a[2], b[6]);
and	(pp[71], a[2], b[7]);
and	(pp[72], a[2], b[8]);
and	(pp[73], a[2], b[9]);
and	(pp[74], a[2], b[10]);
and	(pp[75], a[2], b[11]);
and	(pp[76], a[2], b[12]);
and	(pp[77], a[2], b[13]);
and	(pp[78], a[2], b[14]);
and	(pp[79], a[2], b[15]);
and	(pp[80], a[2], b[16]);
and	(pp[81], a[2], b[17]);
and	(pp[82], a[2], b[18]);
and	(pp[83], a[2], b[19]);
and	(pp[84], a[2], b[20]);
and	(pp[85], a[2], b[21]);
and	(pp[86], a[2], b[22]);
and	(pp[87], a[2], b[23]);
and	(pp[88], a[2], b[24]);
and	(pp[89], a[2], b[25]);
and	(pp[90], a[2], b[26]);
and	(pp[91], a[2], b[27]);
and	(pp[92], a[2], b[28]);
and	(pp[93], a[2], b[29]);
and	(pp[94], a[2], b[30]);
and	(pp[95], a[2], b[31]);
and	(pp[96], a[3], b[0]);
and	(pp[97], a[3], b[1]);
and	(pp[98], a[3], b[2]);
and	(pp[99], a[3], b[3]);
and	(pp[100], a[3], b[4]);
and	(pp[101], a[3], b[5]);
and	(pp[102], a[3], b[6]);
and	(pp[103], a[3], b[7]);
and	(pp[104], a[3], b[8]);
and	(pp[105], a[3], b[9]);
and	(pp[106], a[3], b[10]);
and	(pp[107], a[3], b[11]);
and	(pp[108], a[3], b[12]);
and	(pp[109], a[3], b[13]);
and	(pp[110], a[3], b[14]);
and	(pp[111], a[3], b[15]);
and	(pp[112], a[3], b[16]);
and	(pp[113], a[3], b[17]);
and	(pp[114], a[3], b[18]);
and	(pp[115], a[3], b[19]);
and	(pp[116], a[3], b[20]);
and	(pp[117], a[3], b[21]);
and	(pp[118], a[3], b[22]);
and	(pp[119], a[3], b[23]);
and	(pp[120], a[3], b[24]);
and	(pp[121], a[3], b[25]);
and	(pp[122], a[3], b[26]);
and	(pp[123], a[3], b[27]);
and	(pp[124], a[3], b[28]);
and	(pp[125], a[3], b[29]);
and	(pp[126], a[3], b[30]);
and	(pp[127], a[3], b[31]);
and	(pp[128], a[4], b[0]);
and	(pp[129], a[4], b[1]);
and	(pp[130], a[4], b[2]);
and	(pp[131], a[4], b[3]);
and	(pp[132], a[4], b[4]);
and	(pp[133], a[4], b[5]);
and	(pp[134], a[4], b[6]);
and	(pp[135], a[4], b[7]);
and	(pp[136], a[4], b[8]);
and	(pp[137], a[4], b[9]);
and	(pp[138], a[4], b[10]);
and	(pp[139], a[4], b[11]);
and	(pp[140], a[4], b[12]);
and	(pp[141], a[4], b[13]);
and	(pp[142], a[4], b[14]);
and	(pp[143], a[4], b[15]);
and	(pp[144], a[4], b[16]);
and	(pp[145], a[4], b[17]);
and	(pp[146], a[4], b[18]);
and	(pp[147], a[4], b[19]);
and	(pp[148], a[4], b[20]);
and	(pp[149], a[4], b[21]);
and	(pp[150], a[4], b[22]);
and	(pp[151], a[4], b[23]);
and	(pp[152], a[4], b[24]);
and	(pp[153], a[4], b[25]);
and	(pp[154], a[4], b[26]);
and	(pp[155], a[4], b[27]);
and	(pp[156], a[4], b[28]);
and	(pp[157], a[4], b[29]);
and	(pp[158], a[4], b[30]);
and	(pp[159], a[4], b[31]);
and	(pp[160], a[5], b[0]);
and	(pp[161], a[5], b[1]);
and	(pp[162], a[5], b[2]);
and	(pp[163], a[5], b[3]);
and	(pp[164], a[5], b[4]);
and	(pp[165], a[5], b[5]);
and	(pp[166], a[5], b[6]);
and	(pp[167], a[5], b[7]);
and	(pp[168], a[5], b[8]);
and	(pp[169], a[5], b[9]);
and	(pp[170], a[5], b[10]);
and	(pp[171], a[5], b[11]);
and	(pp[172], a[5], b[12]);
and	(pp[173], a[5], b[13]);
and	(pp[174], a[5], b[14]);
and	(pp[175], a[5], b[15]);
and	(pp[176], a[5], b[16]);
and	(pp[177], a[5], b[17]);
and	(pp[178], a[5], b[18]);
and	(pp[179], a[5], b[19]);
and	(pp[180], a[5], b[20]);
and	(pp[181], a[5], b[21]);
and	(pp[182], a[5], b[22]);
and	(pp[183], a[5], b[23]);
and	(pp[184], a[5], b[24]);
and	(pp[185], a[5], b[25]);
and	(pp[186], a[5], b[26]);
and	(pp[187], a[5], b[27]);
and	(pp[188], a[5], b[28]);
and	(pp[189], a[5], b[29]);
and	(pp[190], a[5], b[30]);
and	(pp[191], a[5], b[31]);
and	(pp[192], a[6], b[0]);
and	(pp[193], a[6], b[1]);
and	(pp[194], a[6], b[2]);
and	(pp[195], a[6], b[3]);
and	(pp[196], a[6], b[4]);
and	(pp[197], a[6], b[5]);
and	(pp[198], a[6], b[6]);
and	(pp[199], a[6], b[7]);
and	(pp[200], a[6], b[8]);
and	(pp[201], a[6], b[9]);
and	(pp[202], a[6], b[10]);
and	(pp[203], a[6], b[11]);
and	(pp[204], a[6], b[12]);
and	(pp[205], a[6], b[13]);
and	(pp[206], a[6], b[14]);
and	(pp[207], a[6], b[15]);
and	(pp[208], a[6], b[16]);
and	(pp[209], a[6], b[17]);
and	(pp[210], a[6], b[18]);
and	(pp[211], a[6], b[19]);
and	(pp[212], a[6], b[20]);
and	(pp[213], a[6], b[21]);
and	(pp[214], a[6], b[22]);
and	(pp[215], a[6], b[23]);
and	(pp[216], a[6], b[24]);
and	(pp[217], a[6], b[25]);
and	(pp[218], a[6], b[26]);
and	(pp[219], a[6], b[27]);
and	(pp[220], a[6], b[28]);
and	(pp[221], a[6], b[29]);
and	(pp[222], a[6], b[30]);
and	(pp[223], a[6], b[31]);
and	(pp[224], a[7], b[0]);
and	(pp[225], a[7], b[1]);
and	(pp[226], a[7], b[2]);
and	(pp[227], a[7], b[3]);
and	(pp[228], a[7], b[4]);
and	(pp[229], a[7], b[5]);
and	(pp[230], a[7], b[6]);
and	(pp[231], a[7], b[7]);
and	(pp[232], a[7], b[8]);
and	(pp[233], a[7], b[9]);
and	(pp[234], a[7], b[10]);
and	(pp[235], a[7], b[11]);
and	(pp[236], a[7], b[12]);
and	(pp[237], a[7], b[13]);
and	(pp[238], a[7], b[14]);
and	(pp[239], a[7], b[15]);
and	(pp[240], a[7], b[16]);
and	(pp[241], a[7], b[17]);
and	(pp[242], a[7], b[18]);
and	(pp[243], a[7], b[19]);
and	(pp[244], a[7], b[20]);
and	(pp[245], a[7], b[21]);
and	(pp[246], a[7], b[22]);
and	(pp[247], a[7], b[23]);
and	(pp[248], a[7], b[24]);
and	(pp[249], a[7], b[25]);
and	(pp[250], a[7], b[26]);
and	(pp[251], a[7], b[27]);
and	(pp[252], a[7], b[28]);
and	(pp[253], a[7], b[29]);
and	(pp[254], a[7], b[30]);
and	(pp[255], a[7], b[31]);
and	(pp[256], a[8], b[0]);
and	(pp[257], a[8], b[1]);
and	(pp[258], a[8], b[2]);
and	(pp[259], a[8], b[3]);
and	(pp[260], a[8], b[4]);
and	(pp[261], a[8], b[5]);
and	(pp[262], a[8], b[6]);
and	(pp[263], a[8], b[7]);
and	(pp[264], a[8], b[8]);
and	(pp[265], a[8], b[9]);
and	(pp[266], a[8], b[10]);
and	(pp[267], a[8], b[11]);
and	(pp[268], a[8], b[12]);
and	(pp[269], a[8], b[13]);
and	(pp[270], a[8], b[14]);
and	(pp[271], a[8], b[15]);
and	(pp[272], a[8], b[16]);
and	(pp[273], a[8], b[17]);
and	(pp[274], a[8], b[18]);
and	(pp[275], a[8], b[19]);
and	(pp[276], a[8], b[20]);
and	(pp[277], a[8], b[21]);
and	(pp[278], a[8], b[22]);
and	(pp[279], a[8], b[23]);
and	(pp[280], a[8], b[24]);
and	(pp[281], a[8], b[25]);
and	(pp[282], a[8], b[26]);
and	(pp[283], a[8], b[27]);
and	(pp[284], a[8], b[28]);
and	(pp[285], a[8], b[29]);
and	(pp[286], a[8], b[30]);
and	(pp[287], a[8], b[31]);
and	(pp[288], a[9], b[0]);
and	(pp[289], a[9], b[1]);
and	(pp[290], a[9], b[2]);
and	(pp[291], a[9], b[3]);
and	(pp[292], a[9], b[4]);
and	(pp[293], a[9], b[5]);
and	(pp[294], a[9], b[6]);
and	(pp[295], a[9], b[7]);
and	(pp[296], a[9], b[8]);
and	(pp[297], a[9], b[9]);
and	(pp[298], a[9], b[10]);
and	(pp[299], a[9], b[11]);
and	(pp[300], a[9], b[12]);
and	(pp[301], a[9], b[13]);
and	(pp[302], a[9], b[14]);
and	(pp[303], a[9], b[15]);
and	(pp[304], a[9], b[16]);
and	(pp[305], a[9], b[17]);
and	(pp[306], a[9], b[18]);
and	(pp[307], a[9], b[19]);
and	(pp[308], a[9], b[20]);
and	(pp[309], a[9], b[21]);
and	(pp[310], a[9], b[22]);
and	(pp[311], a[9], b[23]);
and	(pp[312], a[9], b[24]);
and	(pp[313], a[9], b[25]);
and	(pp[314], a[9], b[26]);
and	(pp[315], a[9], b[27]);
and	(pp[316], a[9], b[28]);
and	(pp[317], a[9], b[29]);
and	(pp[318], a[9], b[30]);
and	(pp[319], a[9], b[31]);
and	(pp[320], a[10], b[0]);
and	(pp[321], a[10], b[1]);
and	(pp[322], a[10], b[2]);
and	(pp[323], a[10], b[3]);
and	(pp[324], a[10], b[4]);
and	(pp[325], a[10], b[5]);
and	(pp[326], a[10], b[6]);
and	(pp[327], a[10], b[7]);
and	(pp[328], a[10], b[8]);
and	(pp[329], a[10], b[9]);
and	(pp[330], a[10], b[10]);
and	(pp[331], a[10], b[11]);
and	(pp[332], a[10], b[12]);
and	(pp[333], a[10], b[13]);
and	(pp[334], a[10], b[14]);
and	(pp[335], a[10], b[15]);
and	(pp[336], a[10], b[16]);
and	(pp[337], a[10], b[17]);
and	(pp[338], a[10], b[18]);
and	(pp[339], a[10], b[19]);
and	(pp[340], a[10], b[20]);
and	(pp[341], a[10], b[21]);
and	(pp[342], a[10], b[22]);
and	(pp[343], a[10], b[23]);
and	(pp[344], a[10], b[24]);
and	(pp[345], a[10], b[25]);
and	(pp[346], a[10], b[26]);
and	(pp[347], a[10], b[27]);
and	(pp[348], a[10], b[28]);
and	(pp[349], a[10], b[29]);
and	(pp[350], a[10], b[30]);
and	(pp[351], a[10], b[31]);
and	(pp[352], a[11], b[0]);
and	(pp[353], a[11], b[1]);
and	(pp[354], a[11], b[2]);
and	(pp[355], a[11], b[3]);
and	(pp[356], a[11], b[4]);
and	(pp[357], a[11], b[5]);
and	(pp[358], a[11], b[6]);
and	(pp[359], a[11], b[7]);
and	(pp[360], a[11], b[8]);
and	(pp[361], a[11], b[9]);
and	(pp[362], a[11], b[10]);
and	(pp[363], a[11], b[11]);
and	(pp[364], a[11], b[12]);
and	(pp[365], a[11], b[13]);
and	(pp[366], a[11], b[14]);
and	(pp[367], a[11], b[15]);
and	(pp[368], a[11], b[16]);
and	(pp[369], a[11], b[17]);
and	(pp[370], a[11], b[18]);
and	(pp[371], a[11], b[19]);
and	(pp[372], a[11], b[20]);
and	(pp[373], a[11], b[21]);
and	(pp[374], a[11], b[22]);
and	(pp[375], a[11], b[23]);
and	(pp[376], a[11], b[24]);
and	(pp[377], a[11], b[25]);
and	(pp[378], a[11], b[26]);
and	(pp[379], a[11], b[27]);
and	(pp[380], a[11], b[28]);
and	(pp[381], a[11], b[29]);
and	(pp[382], a[11], b[30]);
and	(pp[383], a[11], b[31]);
and	(pp[384], a[12], b[0]);
and	(pp[385], a[12], b[1]);
and	(pp[386], a[12], b[2]);
and	(pp[387], a[12], b[3]);
and	(pp[388], a[12], b[4]);
and	(pp[389], a[12], b[5]);
and	(pp[390], a[12], b[6]);
and	(pp[391], a[12], b[7]);
and	(pp[392], a[12], b[8]);
and	(pp[393], a[12], b[9]);
and	(pp[394], a[12], b[10]);
and	(pp[395], a[12], b[11]);
and	(pp[396], a[12], b[12]);
and	(pp[397], a[12], b[13]);
and	(pp[398], a[12], b[14]);
and	(pp[399], a[12], b[15]);
and	(pp[400], a[12], b[16]);
and	(pp[401], a[12], b[17]);
and	(pp[402], a[12], b[18]);
and	(pp[403], a[12], b[19]);
and	(pp[404], a[12], b[20]);
and	(pp[405], a[12], b[21]);
and	(pp[406], a[12], b[22]);
and	(pp[407], a[12], b[23]);
and	(pp[408], a[12], b[24]);
and	(pp[409], a[12], b[25]);
and	(pp[410], a[12], b[26]);
and	(pp[411], a[12], b[27]);
and	(pp[412], a[12], b[28]);
and	(pp[413], a[12], b[29]);
and	(pp[414], a[12], b[30]);
and	(pp[415], a[12], b[31]);
and	(pp[416], a[13], b[0]);
and	(pp[417], a[13], b[1]);
and	(pp[418], a[13], b[2]);
and	(pp[419], a[13], b[3]);
and	(pp[420], a[13], b[4]);
and	(pp[421], a[13], b[5]);
and	(pp[422], a[13], b[6]);
and	(pp[423], a[13], b[7]);
and	(pp[424], a[13], b[8]);
and	(pp[425], a[13], b[9]);
and	(pp[426], a[13], b[10]);
and	(pp[427], a[13], b[11]);
and	(pp[428], a[13], b[12]);
and	(pp[429], a[13], b[13]);
and	(pp[430], a[13], b[14]);
and	(pp[431], a[13], b[15]);
and	(pp[432], a[13], b[16]);
and	(pp[433], a[13], b[17]);
and	(pp[434], a[13], b[18]);
and	(pp[435], a[13], b[19]);
and	(pp[436], a[13], b[20]);
and	(pp[437], a[13], b[21]);
and	(pp[438], a[13], b[22]);
and	(pp[439], a[13], b[23]);
and	(pp[440], a[13], b[24]);
and	(pp[441], a[13], b[25]);
and	(pp[442], a[13], b[26]);
and	(pp[443], a[13], b[27]);
and	(pp[444], a[13], b[28]);
and	(pp[445], a[13], b[29]);
and	(pp[446], a[13], b[30]);
and	(pp[447], a[13], b[31]);
and	(pp[448], a[14], b[0]);
and	(pp[449], a[14], b[1]);
and	(pp[450], a[14], b[2]);
and	(pp[451], a[14], b[3]);
and	(pp[452], a[14], b[4]);
and	(pp[453], a[14], b[5]);
and	(pp[454], a[14], b[6]);
and	(pp[455], a[14], b[7]);
and	(pp[456], a[14], b[8]);
and	(pp[457], a[14], b[9]);
and	(pp[458], a[14], b[10]);
and	(pp[459], a[14], b[11]);
and	(pp[460], a[14], b[12]);
and	(pp[461], a[14], b[13]);
and	(pp[462], a[14], b[14]);
and	(pp[463], a[14], b[15]);
and	(pp[464], a[14], b[16]);
and	(pp[465], a[14], b[17]);
and	(pp[466], a[14], b[18]);
and	(pp[467], a[14], b[19]);
and	(pp[468], a[14], b[20]);
and	(pp[469], a[14], b[21]);
and	(pp[470], a[14], b[22]);
and	(pp[471], a[14], b[23]);
and	(pp[472], a[14], b[24]);
and	(pp[473], a[14], b[25]);
and	(pp[474], a[14], b[26]);
and	(pp[475], a[14], b[27]);
and	(pp[476], a[14], b[28]);
and	(pp[477], a[14], b[29]);
and	(pp[478], a[14], b[30]);
and	(pp[479], a[14], b[31]);
and	(pp[480], a[15], b[0]);
and	(pp[481], a[15], b[1]);
and	(pp[482], a[15], b[2]);
and	(pp[483], a[15], b[3]);
and	(pp[484], a[15], b[4]);
and	(pp[485], a[15], b[5]);
and	(pp[486], a[15], b[6]);
and	(pp[487], a[15], b[7]);
and	(pp[488], a[15], b[8]);
and	(pp[489], a[15], b[9]);
and	(pp[490], a[15], b[10]);
and	(pp[491], a[15], b[11]);
and	(pp[492], a[15], b[12]);
and	(pp[493], a[15], b[13]);
and	(pp[494], a[15], b[14]);
and	(pp[495], a[15], b[15]);
and	(pp[496], a[15], b[16]);
and	(pp[497], a[15], b[17]);
and	(pp[498], a[15], b[18]);
and	(pp[499], a[15], b[19]);
and	(pp[500], a[15], b[20]);
and	(pp[501], a[15], b[21]);
and	(pp[502], a[15], b[22]);
and	(pp[503], a[15], b[23]);
and	(pp[504], a[15], b[24]);
and	(pp[505], a[15], b[25]);
and	(pp[506], a[15], b[26]);
and	(pp[507], a[15], b[27]);
and	(pp[508], a[15], b[28]);
and	(pp[509], a[15], b[29]);
and	(pp[510], a[15], b[30]);
and	(pp[511], a[15], b[31]);
and	(pp[512], a[16], b[0]);
and	(pp[513], a[16], b[1]);
and	(pp[514], a[16], b[2]);
and	(pp[515], a[16], b[3]);
and	(pp[516], a[16], b[4]);
and	(pp[517], a[16], b[5]);
and	(pp[518], a[16], b[6]);
and	(pp[519], a[16], b[7]);
and	(pp[520], a[16], b[8]);
and	(pp[521], a[16], b[9]);
and	(pp[522], a[16], b[10]);
and	(pp[523], a[16], b[11]);
and	(pp[524], a[16], b[12]);
and	(pp[525], a[16], b[13]);
and	(pp[526], a[16], b[14]);
and	(pp[527], a[16], b[15]);
and	(pp[528], a[16], b[16]);
and	(pp[529], a[16], b[17]);
and	(pp[530], a[16], b[18]);
and	(pp[531], a[16], b[19]);
and	(pp[532], a[16], b[20]);
and	(pp[533], a[16], b[21]);
and	(pp[534], a[16], b[22]);
and	(pp[535], a[16], b[23]);
and	(pp[536], a[16], b[24]);
and	(pp[537], a[16], b[25]);
and	(pp[538], a[16], b[26]);
and	(pp[539], a[16], b[27]);
and	(pp[540], a[16], b[28]);
and	(pp[541], a[16], b[29]);
and	(pp[542], a[16], b[30]);
and	(pp[543], a[16], b[31]);
and	(pp[544], a[17], b[0]);
and	(pp[545], a[17], b[1]);
and	(pp[546], a[17], b[2]);
and	(pp[547], a[17], b[3]);
and	(pp[548], a[17], b[4]);
and	(pp[549], a[17], b[5]);
and	(pp[550], a[17], b[6]);
and	(pp[551], a[17], b[7]);
and	(pp[552], a[17], b[8]);
and	(pp[553], a[17], b[9]);
and	(pp[554], a[17], b[10]);
and	(pp[555], a[17], b[11]);
and	(pp[556], a[17], b[12]);
and	(pp[557], a[17], b[13]);
and	(pp[558], a[17], b[14]);
and	(pp[559], a[17], b[15]);
and	(pp[560], a[17], b[16]);
and	(pp[561], a[17], b[17]);
and	(pp[562], a[17], b[18]);
and	(pp[563], a[17], b[19]);
and	(pp[564], a[17], b[20]);
and	(pp[565], a[17], b[21]);
and	(pp[566], a[17], b[22]);
and	(pp[567], a[17], b[23]);
and	(pp[568], a[17], b[24]);
and	(pp[569], a[17], b[25]);
and	(pp[570], a[17], b[26]);
and	(pp[571], a[17], b[27]);
and	(pp[572], a[17], b[28]);
and	(pp[573], a[17], b[29]);
and	(pp[574], a[17], b[30]);
and	(pp[575], a[17], b[31]);
and	(pp[576], a[18], b[0]);
and	(pp[577], a[18], b[1]);
and	(pp[578], a[18], b[2]);
and	(pp[579], a[18], b[3]);
and	(pp[580], a[18], b[4]);
and	(pp[581], a[18], b[5]);
and	(pp[582], a[18], b[6]);
and	(pp[583], a[18], b[7]);
and	(pp[584], a[18], b[8]);
and	(pp[585], a[18], b[9]);
and	(pp[586], a[18], b[10]);
and	(pp[587], a[18], b[11]);
and	(pp[588], a[18], b[12]);
and	(pp[589], a[18], b[13]);
and	(pp[590], a[18], b[14]);
and	(pp[591], a[18], b[15]);
and	(pp[592], a[18], b[16]);
and	(pp[593], a[18], b[17]);
and	(pp[594], a[18], b[18]);
and	(pp[595], a[18], b[19]);
and	(pp[596], a[18], b[20]);
and	(pp[597], a[18], b[21]);
and	(pp[598], a[18], b[22]);
and	(pp[599], a[18], b[23]);
and	(pp[600], a[18], b[24]);
and	(pp[601], a[18], b[25]);
and	(pp[602], a[18], b[26]);
and	(pp[603], a[18], b[27]);
and	(pp[604], a[18], b[28]);
and	(pp[605], a[18], b[29]);
and	(pp[606], a[18], b[30]);
and	(pp[607], a[18], b[31]);
and	(pp[608], a[19], b[0]);
and	(pp[609], a[19], b[1]);
and	(pp[610], a[19], b[2]);
and	(pp[611], a[19], b[3]);
and	(pp[612], a[19], b[4]);
and	(pp[613], a[19], b[5]);
and	(pp[614], a[19], b[6]);
and	(pp[615], a[19], b[7]);
and	(pp[616], a[19], b[8]);
and	(pp[617], a[19], b[9]);
and	(pp[618], a[19], b[10]);
and	(pp[619], a[19], b[11]);
and	(pp[620], a[19], b[12]);
and	(pp[621], a[19], b[13]);
and	(pp[622], a[19], b[14]);
and	(pp[623], a[19], b[15]);
and	(pp[624], a[19], b[16]);
and	(pp[625], a[19], b[17]);
and	(pp[626], a[19], b[18]);
and	(pp[627], a[19], b[19]);
and	(pp[628], a[19], b[20]);
and	(pp[629], a[19], b[21]);
and	(pp[630], a[19], b[22]);
and	(pp[631], a[19], b[23]);
and	(pp[632], a[19], b[24]);
and	(pp[633], a[19], b[25]);
and	(pp[634], a[19], b[26]);
and	(pp[635], a[19], b[27]);
and	(pp[636], a[19], b[28]);
and	(pp[637], a[19], b[29]);
and	(pp[638], a[19], b[30]);
and	(pp[639], a[19], b[31]);
and	(pp[640], a[20], b[0]);
and	(pp[641], a[20], b[1]);
and	(pp[642], a[20], b[2]);
and	(pp[643], a[20], b[3]);
and	(pp[644], a[20], b[4]);
and	(pp[645], a[20], b[5]);
and	(pp[646], a[20], b[6]);
and	(pp[647], a[20], b[7]);
and	(pp[648], a[20], b[8]);
and	(pp[649], a[20], b[9]);
and	(pp[650], a[20], b[10]);
and	(pp[651], a[20], b[11]);
and	(pp[652], a[20], b[12]);
and	(pp[653], a[20], b[13]);
and	(pp[654], a[20], b[14]);
and	(pp[655], a[20], b[15]);
and	(pp[656], a[20], b[16]);
and	(pp[657], a[20], b[17]);
and	(pp[658], a[20], b[18]);
and	(pp[659], a[20], b[19]);
and	(pp[660], a[20], b[20]);
and	(pp[661], a[20], b[21]);
and	(pp[662], a[20], b[22]);
and	(pp[663], a[20], b[23]);
and	(pp[664], a[20], b[24]);
and	(pp[665], a[20], b[25]);
and	(pp[666], a[20], b[26]);
and	(pp[667], a[20], b[27]);
and	(pp[668], a[20], b[28]);
and	(pp[669], a[20], b[29]);
and	(pp[670], a[20], b[30]);
and	(pp[671], a[20], b[31]);
and	(pp[672], a[21], b[0]);
and	(pp[673], a[21], b[1]);
and	(pp[674], a[21], b[2]);
and	(pp[675], a[21], b[3]);
and	(pp[676], a[21], b[4]);
and	(pp[677], a[21], b[5]);
and	(pp[678], a[21], b[6]);
and	(pp[679], a[21], b[7]);
and	(pp[680], a[21], b[8]);
and	(pp[681], a[21], b[9]);
and	(pp[682], a[21], b[10]);
and	(pp[683], a[21], b[11]);
and	(pp[684], a[21], b[12]);
and	(pp[685], a[21], b[13]);
and	(pp[686], a[21], b[14]);
and	(pp[687], a[21], b[15]);
and	(pp[688], a[21], b[16]);
and	(pp[689], a[21], b[17]);
and	(pp[690], a[21], b[18]);
and	(pp[691], a[21], b[19]);
and	(pp[692], a[21], b[20]);
and	(pp[693], a[21], b[21]);
and	(pp[694], a[21], b[22]);
and	(pp[695], a[21], b[23]);
and	(pp[696], a[21], b[24]);
and	(pp[697], a[21], b[25]);
and	(pp[698], a[21], b[26]);
and	(pp[699], a[21], b[27]);
and	(pp[700], a[21], b[28]);
and	(pp[701], a[21], b[29]);
and	(pp[702], a[21], b[30]);
and	(pp[703], a[21], b[31]);
and	(pp[704], a[22], b[0]);
and	(pp[705], a[22], b[1]);
and	(pp[706], a[22], b[2]);
and	(pp[707], a[22], b[3]);
and	(pp[708], a[22], b[4]);
and	(pp[709], a[22], b[5]);
and	(pp[710], a[22], b[6]);
and	(pp[711], a[22], b[7]);
and	(pp[712], a[22], b[8]);
and	(pp[713], a[22], b[9]);
and	(pp[714], a[22], b[10]);
and	(pp[715], a[22], b[11]);
and	(pp[716], a[22], b[12]);
and	(pp[717], a[22], b[13]);
and	(pp[718], a[22], b[14]);
and	(pp[719], a[22], b[15]);
and	(pp[720], a[22], b[16]);
and	(pp[721], a[22], b[17]);
and	(pp[722], a[22], b[18]);
and	(pp[723], a[22], b[19]);
and	(pp[724], a[22], b[20]);
and	(pp[725], a[22], b[21]);
and	(pp[726], a[22], b[22]);
and	(pp[727], a[22], b[23]);
and	(pp[728], a[22], b[24]);
and	(pp[729], a[22], b[25]);
and	(pp[730], a[22], b[26]);
and	(pp[731], a[22], b[27]);
and	(pp[732], a[22], b[28]);
and	(pp[733], a[22], b[29]);
and	(pp[734], a[22], b[30]);
and	(pp[735], a[22], b[31]);
and	(pp[736], a[23], b[0]);
and	(pp[737], a[23], b[1]);
and	(pp[738], a[23], b[2]);
and	(pp[739], a[23], b[3]);
and	(pp[740], a[23], b[4]);
and	(pp[741], a[23], b[5]);
and	(pp[742], a[23], b[6]);
and	(pp[743], a[23], b[7]);
and	(pp[744], a[23], b[8]);
and	(pp[745], a[23], b[9]);
and	(pp[746], a[23], b[10]);
and	(pp[747], a[23], b[11]);
and	(pp[748], a[23], b[12]);
and	(pp[749], a[23], b[13]);
and	(pp[750], a[23], b[14]);
and	(pp[751], a[23], b[15]);
and	(pp[752], a[23], b[16]);
and	(pp[753], a[23], b[17]);
and	(pp[754], a[23], b[18]);
and	(pp[755], a[23], b[19]);
and	(pp[756], a[23], b[20]);
and	(pp[757], a[23], b[21]);
and	(pp[758], a[23], b[22]);
and	(pp[759], a[23], b[23]);
and	(pp[760], a[23], b[24]);
and	(pp[761], a[23], b[25]);
and	(pp[762], a[23], b[26]);
and	(pp[763], a[23], b[27]);
and	(pp[764], a[23], b[28]);
and	(pp[765], a[23], b[29]);
and	(pp[766], a[23], b[30]);
and	(pp[767], a[23], b[31]);
and	(pp[768], a[24], b[0]);
and	(pp[769], a[24], b[1]);
and	(pp[770], a[24], b[2]);
and	(pp[771], a[24], b[3]);
and	(pp[772], a[24], b[4]);
and	(pp[773], a[24], b[5]);
and	(pp[774], a[24], b[6]);
and	(pp[775], a[24], b[7]);
and	(pp[776], a[24], b[8]);
and	(pp[777], a[24], b[9]);
and	(pp[778], a[24], b[10]);
and	(pp[779], a[24], b[11]);
and	(pp[780], a[24], b[12]);
and	(pp[781], a[24], b[13]);
and	(pp[782], a[24], b[14]);
and	(pp[783], a[24], b[15]);
and	(pp[784], a[24], b[16]);
and	(pp[785], a[24], b[17]);
and	(pp[786], a[24], b[18]);
and	(pp[787], a[24], b[19]);
and	(pp[788], a[24], b[20]);
and	(pp[789], a[24], b[21]);
and	(pp[790], a[24], b[22]);
and	(pp[791], a[24], b[23]);
and	(pp[792], a[24], b[24]);
and	(pp[793], a[24], b[25]);
and	(pp[794], a[24], b[26]);
and	(pp[795], a[24], b[27]);
and	(pp[796], a[24], b[28]);
and	(pp[797], a[24], b[29]);
and	(pp[798], a[24], b[30]);
and	(pp[799], a[24], b[31]);
and	(pp[800], a[25], b[0]);
and	(pp[801], a[25], b[1]);
and	(pp[802], a[25], b[2]);
and	(pp[803], a[25], b[3]);
and	(pp[804], a[25], b[4]);
and	(pp[805], a[25], b[5]);
and	(pp[806], a[25], b[6]);
and	(pp[807], a[25], b[7]);
and	(pp[808], a[25], b[8]);
and	(pp[809], a[25], b[9]);
and	(pp[810], a[25], b[10]);
and	(pp[811], a[25], b[11]);
and	(pp[812], a[25], b[12]);
and	(pp[813], a[25], b[13]);
and	(pp[814], a[25], b[14]);
and	(pp[815], a[25], b[15]);
and	(pp[816], a[25], b[16]);
and	(pp[817], a[25], b[17]);
and	(pp[818], a[25], b[18]);
and	(pp[819], a[25], b[19]);
and	(pp[820], a[25], b[20]);
and	(pp[821], a[25], b[21]);
and	(pp[822], a[25], b[22]);
and	(pp[823], a[25], b[23]);
and	(pp[824], a[25], b[24]);
and	(pp[825], a[25], b[25]);
and	(pp[826], a[25], b[26]);
and	(pp[827], a[25], b[27]);
and	(pp[828], a[25], b[28]);
and	(pp[829], a[25], b[29]);
and	(pp[830], a[25], b[30]);
and	(pp[831], a[25], b[31]);
and	(pp[832], a[26], b[0]);
and	(pp[833], a[26], b[1]);
and	(pp[834], a[26], b[2]);
and	(pp[835], a[26], b[3]);
and	(pp[836], a[26], b[4]);
and	(pp[837], a[26], b[5]);
and	(pp[838], a[26], b[6]);
and	(pp[839], a[26], b[7]);
and	(pp[840], a[26], b[8]);
and	(pp[841], a[26], b[9]);
and	(pp[842], a[26], b[10]);
and	(pp[843], a[26], b[11]);
and	(pp[844], a[26], b[12]);
and	(pp[845], a[26], b[13]);
and	(pp[846], a[26], b[14]);
and	(pp[847], a[26], b[15]);
and	(pp[848], a[26], b[16]);
and	(pp[849], a[26], b[17]);
and	(pp[850], a[26], b[18]);
and	(pp[851], a[26], b[19]);
and	(pp[852], a[26], b[20]);
and	(pp[853], a[26], b[21]);
and	(pp[854], a[26], b[22]);
and	(pp[855], a[26], b[23]);
and	(pp[856], a[26], b[24]);
and	(pp[857], a[26], b[25]);
and	(pp[858], a[26], b[26]);
and	(pp[859], a[26], b[27]);
and	(pp[860], a[26], b[28]);
and	(pp[861], a[26], b[29]);
and	(pp[862], a[26], b[30]);
and	(pp[863], a[26], b[31]);
and	(pp[864], a[27], b[0]);
and	(pp[865], a[27], b[1]);
and	(pp[866], a[27], b[2]);
and	(pp[867], a[27], b[3]);
and	(pp[868], a[27], b[4]);
and	(pp[869], a[27], b[5]);
and	(pp[870], a[27], b[6]);
and	(pp[871], a[27], b[7]);
and	(pp[872], a[27], b[8]);
and	(pp[873], a[27], b[9]);
and	(pp[874], a[27], b[10]);
and	(pp[875], a[27], b[11]);
and	(pp[876], a[27], b[12]);
and	(pp[877], a[27], b[13]);
and	(pp[878], a[27], b[14]);
and	(pp[879], a[27], b[15]);
and	(pp[880], a[27], b[16]);
and	(pp[881], a[27], b[17]);
and	(pp[882], a[27], b[18]);
and	(pp[883], a[27], b[19]);
and	(pp[884], a[27], b[20]);
and	(pp[885], a[27], b[21]);
and	(pp[886], a[27], b[22]);
and	(pp[887], a[27], b[23]);
and	(pp[888], a[27], b[24]);
and	(pp[889], a[27], b[25]);
and	(pp[890], a[27], b[26]);
and	(pp[891], a[27], b[27]);
and	(pp[892], a[27], b[28]);
and	(pp[893], a[27], b[29]);
and	(pp[894], a[27], b[30]);
and	(pp[895], a[27], b[31]);
and	(pp[896], a[28], b[0]);
and	(pp[897], a[28], b[1]);
and	(pp[898], a[28], b[2]);
and	(pp[899], a[28], b[3]);
and	(pp[900], a[28], b[4]);
and	(pp[901], a[28], b[5]);
and	(pp[902], a[28], b[6]);
and	(pp[903], a[28], b[7]);
and	(pp[904], a[28], b[8]);
and	(pp[905], a[28], b[9]);
and	(pp[906], a[28], b[10]);
and	(pp[907], a[28], b[11]);
and	(pp[908], a[28], b[12]);
and	(pp[909], a[28], b[13]);
and	(pp[910], a[28], b[14]);
and	(pp[911], a[28], b[15]);
and	(pp[912], a[28], b[16]);
and	(pp[913], a[28], b[17]);
and	(pp[914], a[28], b[18]);
and	(pp[915], a[28], b[19]);
and	(pp[916], a[28], b[20]);
and	(pp[917], a[28], b[21]);
and	(pp[918], a[28], b[22]);
and	(pp[919], a[28], b[23]);
and	(pp[920], a[28], b[24]);
and	(pp[921], a[28], b[25]);
and	(pp[922], a[28], b[26]);
and	(pp[923], a[28], b[27]);
and	(pp[924], a[28], b[28]);
and	(pp[925], a[28], b[29]);
and	(pp[926], a[28], b[30]);
and	(pp[927], a[28], b[31]);
and	(pp[928], a[29], b[0]);
and	(pp[929], a[29], b[1]);
and	(pp[930], a[29], b[2]);
and	(pp[931], a[29], b[3]);
and	(pp[932], a[29], b[4]);
and	(pp[933], a[29], b[5]);
and	(pp[934], a[29], b[6]);
and	(pp[935], a[29], b[7]);
and	(pp[936], a[29], b[8]);
and	(pp[937], a[29], b[9]);
and	(pp[938], a[29], b[10]);
and	(pp[939], a[29], b[11]);
and	(pp[940], a[29], b[12]);
and	(pp[941], a[29], b[13]);
and	(pp[942], a[29], b[14]);
and	(pp[943], a[29], b[15]);
and	(pp[944], a[29], b[16]);
and	(pp[945], a[29], b[17]);
and	(pp[946], a[29], b[18]);
and	(pp[947], a[29], b[19]);
and	(pp[948], a[29], b[20]);
and	(pp[949], a[29], b[21]);
and	(pp[950], a[29], b[22]);
and	(pp[951], a[29], b[23]);
and	(pp[952], a[29], b[24]);
and	(pp[953], a[29], b[25]);
and	(pp[954], a[29], b[26]);
and	(pp[955], a[29], b[27]);
and	(pp[956], a[29], b[28]);
and	(pp[957], a[29], b[29]);
and	(pp[958], a[29], b[30]);
and	(pp[959], a[29], b[31]);
and	(pp[960], a[30], b[0]);
and	(pp[961], a[30], b[1]);
and	(pp[962], a[30], b[2]);
and	(pp[963], a[30], b[3]);
and	(pp[964], a[30], b[4]);
and	(pp[965], a[30], b[5]);
and	(pp[966], a[30], b[6]);
and	(pp[967], a[30], b[7]);
and	(pp[968], a[30], b[8]);
and	(pp[969], a[30], b[9]);
and	(pp[970], a[30], b[10]);
and	(pp[971], a[30], b[11]);
and	(pp[972], a[30], b[12]);
and	(pp[973], a[30], b[13]);
and	(pp[974], a[30], b[14]);
and	(pp[975], a[30], b[15]);
and	(pp[976], a[30], b[16]);
and	(pp[977], a[30], b[17]);
and	(pp[978], a[30], b[18]);
and	(pp[979], a[30], b[19]);
and	(pp[980], a[30], b[20]);
and	(pp[981], a[30], b[21]);
and	(pp[982], a[30], b[22]);
and	(pp[983], a[30], b[23]);
and	(pp[984], a[30], b[24]);
and	(pp[985], a[30], b[25]);
and	(pp[986], a[30], b[26]);
and	(pp[987], a[30], b[27]);
and	(pp[988], a[30], b[28]);
and	(pp[989], a[30], b[29]);
and	(pp[990], a[30], b[30]);
and	(pp[991], a[30], b[31]);
and	(pp[992], a[31], b[0]);
and	(pp[993], a[31], b[1]);
and	(pp[994], a[31], b[2]);
and	(pp[995], a[31], b[3]);
and	(pp[996], a[31], b[4]);
and	(pp[997], a[31], b[5]);
and	(pp[998], a[31], b[6]);
and	(pp[999], a[31], b[7]);
and	(pp[1000], a[31], b[8]);
and	(pp[1001], a[31], b[9]);
and	(pp[1002], a[31], b[10]);
and	(pp[1003], a[31], b[11]);
and	(pp[1004], a[31], b[12]);
and	(pp[1005], a[31], b[13]);
and	(pp[1006], a[31], b[14]);
and	(pp[1007], a[31], b[15]);
and	(pp[1008], a[31], b[16]);
and	(pp[1009], a[31], b[17]);
and	(pp[1010], a[31], b[18]);
and	(pp[1011], a[31], b[19]);
and	(pp[1012], a[31], b[20]);
and	(pp[1013], a[31], b[21]);
and	(pp[1014], a[31], b[22]);
and	(pp[1015], a[31], b[23]);
and	(pp[1016], a[31], b[24]);
and	(pp[1017], a[31], b[25]);
and	(pp[1018], a[31], b[26]);
and	(pp[1019], a[31], b[27]);
and	(pp[1020], a[31], b[28]);
and	(pp[1021], a[31], b[29]);
and	(pp[1022], a[31], b[30]);
and	(pp[1023], a[31], b[31]);
//Posible pipline
always @(posedge clk) begin
	pp_reg <= pp;
	ProcConditon_reg[0] <= PDone_in;
end


HA	inst1025	(pp_reg[32], pp_reg[1], m[1], r1c[0]);
FA	inst1026	(pp_reg[33], pp_reg[2], r1c[0], r1s[1], r1c[1]);
FA	inst1027	(pp_reg[34], pp_reg[3], r1c[1], r1s[2], r1c[2]);
FA	inst1028	(pp_reg[35], pp_reg[4], r1c[2], r1s[3], r1c[3]);
FA	inst1029	(pp_reg[36], pp_reg[5], r1c[3], r1s[4], r1c[4]);
FA	inst1030	(pp_reg[37], pp_reg[6], r1c[4], r1s[5], r1c[5]);
FA	inst1031	(pp_reg[38], pp_reg[7], r1c[5], r1s[6], r1c[6]);
FA	inst1032	(pp_reg[39], pp_reg[8], r1c[6], r1s[7], r1c[7]);
FA	inst1033	(pp_reg[40], pp_reg[9], r1c[7], r1s[8], r1c[8]);
FA	inst1034	(pp_reg[41], pp_reg[10], r1c[8], r1s[9], r1c[9]);
FA	inst1035	(pp_reg[42], pp_reg[11], r1c[9], r1s[10], r1c[10]);
FA	inst1036	(pp_reg[43], pp_reg[12], r1c[10], r1s[11], r1c[11]);
FA	inst1037	(pp_reg[44], pp_reg[13], r1c[11], r1s[12], r1c[12]);
FA	inst1038	(pp_reg[45], pp_reg[14], r1c[12], r1s[13], r1c[13]);
FA	inst1039	(pp_reg[46], pp_reg[15], r1c[13], r1s[14], r1c[14]);
FA	inst1040	(pp_reg[47], pp_reg[16], r1c[14], r1s[15], r1c[15]);
FA	inst1041	(pp_reg[48], pp_reg[17], r1c[15], r1s[16], r1c[16]);
FA	inst1042	(pp_reg[49], pp_reg[18], r1c[16], r1s[17], r1c[17]);
FA	inst1043	(pp_reg[50], pp_reg[19], r1c[17], r1s[18], r1c[18]);
FA	inst1044	(pp_reg[51], pp_reg[20], r1c[18], r1s[19], r1c[19]);
FA	inst1045	(pp_reg[52], pp_reg[21], r1c[19], r1s[20], r1c[20]);
FA	inst1046	(pp_reg[53], pp_reg[22], r1c[20], r1s[21], r1c[21]);
FA	inst1047	(pp_reg[54], pp_reg[23], r1c[21], r1s[22], r1c[22]);
FA	inst1048	(pp_reg[55], pp_reg[24], r1c[22], r1s[23], r1c[23]);
FA	inst1049	(pp_reg[56], pp_reg[25], r1c[23], r1s[24], r1c[24]);
FA	inst1050	(pp_reg[57], pp_reg[26], r1c[24], r1s[25], r1c[25]);
FA	inst1051	(pp_reg[58], pp_reg[27], r1c[25], r1s[26], r1c[26]);
FA	inst1052	(pp_reg[59], pp_reg[28], r1c[26], r1s[27], r1c[27]);
FA	inst1053	(pp_reg[60], pp_reg[29], r1c[27], r1s[28], r1c[28]);
FA	inst1054	(pp_reg[61], pp_reg[30], r1c[28], r1s[29], r1c[29]);
FA	inst1055	(pp_reg[62], pp_reg[31], r1c[29], r1s[30], r1c[30]);
//Posible pipline

always @(posedge clk) begin
	r1s_reg <= r1s;
	rc_last_reg[0] <= r1c[30];
	ProcConditon_reg[1] <= ProcConditon_reg[0];
end

HA	inst1056	(r1s_reg[1], pp_reg[64], m[2], r2c[0]);
FA	inst1057	(r1s_reg[2], pp_reg[65], r2c[0], r2s[1], r2c[1]);
FA	inst1058	(r1s_reg[3], pp_reg[66], r2c[1], r2s[2], r2c[2]);
FA	inst1059	(r1s_reg[4], pp_reg[67], r2c[2], r2s[3], r2c[3]);
FA	inst1060	(r1s_reg[5], pp_reg[68], r2c[3], r2s[4], r2c[4]);
FA	inst1061	(r1s_reg[6], pp_reg[69], r2c[4], r2s[5], r2c[5]);
FA	inst1062	(r1s_reg[7], pp_reg[70], r2c[5], r2s[6], r2c[6]);
FA	inst1063	(r1s_reg[8], pp_reg[71], r2c[6], r2s[7], r2c[7]);
FA	inst1064	(r1s_reg[9], pp_reg[72], r2c[7], r2s[8], r2c[8]);
FA	inst1065	(r1s_reg[10], pp_reg[73], r2c[8], r2s[9], r2c[9]);
FA	inst1066	(r1s_reg[11], pp_reg[74], r2c[9], r2s[10], r2c[10]);
FA	inst1067	(r1s_reg[12], pp_reg[75], r2c[10], r2s[11], r2c[11]);
FA	inst1068	(r1s_reg[13], pp_reg[76], r2c[11], r2s[12], r2c[12]);
FA	inst1069	(r1s_reg[14], pp_reg[77], r2c[12], r2s[13], r2c[13]);
FA	inst1070	(r1s_reg[15], pp_reg[78], r2c[13], r2s[14], r2c[14]);
FA	inst1071	(r1s_reg[16], pp_reg[79], r2c[14], r2s[15], r2c[15]);
FA	inst1072	(r1s_reg[17], pp_reg[80], r2c[15], r2s[16], r2c[16]);
FA	inst1073	(r1s_reg[18], pp_reg[81], r2c[16], r2s[17], r2c[17]);
FA	inst1074	(r1s_reg[19], pp_reg[82], r2c[17], r2s[18], r2c[18]);
FA	inst1075	(r1s_reg[20], pp_reg[83], r2c[18], r2s[19], r2c[19]);
FA	inst1076	(r1s_reg[21], pp_reg[84], r2c[19], r2s[20], r2c[20]);
FA	inst1077	(r1s_reg[22], pp_reg[85], r2c[20], r2s[21], r2c[21]);
FA	inst1078	(r1s_reg[23], pp_reg[86], r2c[21], r2s[22], r2c[22]);
FA	inst1079	(r1s_reg[24], pp_reg[87], r2c[22], r2s[23], r2c[23]);
FA	inst1080	(r1s_reg[25], pp_reg[88], r2c[23], r2s[24], r2c[24]);
FA	inst1081	(r1s_reg[26], pp_reg[89], r2c[24], r2s[25], r2c[25]);
FA	inst1082	(r1s_reg[27], pp_reg[90], r2c[25], r2s[26], r2c[26]);
FA	inst1083	(r1s_reg[28], pp_reg[91], r2c[26], r2s[27], r2c[27]);
FA	inst1084	(r1s_reg[29], pp_reg[92], r2c[27], r2s[28], r2c[28]);
FA	inst1085	(r1s_reg[30], pp_reg[93], r2c[28], r2s[29], r2c[29]);
FA	inst1086	(rc_last_reg[0], pp_reg[63], r2c[29], r2s[30], r2c[30]);
//Posible pipline
always @(posedge clk) begin
	r2s_reg <= r2s;
	rc_last_reg[1] <= r2c[30];
	ProcConditon_reg[2] <= ProcConditon_reg[1];
end

HA	inst1087	(r2s_reg[1], pp_reg[96], m[3], r3c[0]);
FA	inst1088	(r2s_reg[2], pp_reg[97], r3c[0], r3s[1], r3c[1]);
FA	inst1089	(r2s_reg[3], pp_reg[98], r3c[1], r3s[2], r3c[2]);
FA	inst1090	(r2s_reg[4], pp_reg[99], r3c[2], r3s[3], r3c[3]);
FA	inst1091	(r2s_reg[5], pp_reg[100], r3c[3], r3s[4], r3c[4]);
FA	inst1092	(r2s_reg[6], pp_reg[101], r3c[4], r3s[5], r3c[5]);
FA	inst1093	(r2s_reg[7], pp_reg[102], r3c[5], r3s[6], r3c[6]);
FA	inst1094	(r2s_reg[8], pp_reg[103], r3c[6], r3s[7], r3c[7]);
FA	inst1095	(r2s_reg[9], pp_reg[104], r3c[7], r3s[8], r3c[8]);
FA	inst1096	(r2s_reg[10], pp_reg[105], r3c[8], r3s[9], r3c[9]);
FA	inst1097	(r2s_reg[11], pp_reg[106], r3c[9], r3s[10], r3c[10]);
FA	inst1098	(r2s_reg[12], pp_reg[107], r3c[10], r3s[11], r3c[11]);
FA	inst1099	(r2s_reg[13], pp_reg[108], r3c[11], r3s[12], r3c[12]);
FA	inst1100	(r2s_reg[14], pp_reg[109], r3c[12], r3s[13], r3c[13]);
FA	inst1101	(r2s_reg[15], pp_reg[110], r3c[13], r3s[14], r3c[14]);
FA	inst1102	(r2s_reg[16], pp_reg[111], r3c[14], r3s[15], r3c[15]);
FA	inst1103	(r2s_reg[17], pp_reg[112], r3c[15], r3s[16], r3c[16]);
FA	inst1104	(r2s_reg[18], pp_reg[113], r3c[16], r3s[17], r3c[17]);
FA	inst1105	(r2s_reg[19], pp_reg[114], r3c[17], r3s[18], r3c[18]);
FA	inst1106	(r2s_reg[20], pp_reg[115], r3c[18], r3s[19], r3c[19]);
FA	inst1107	(r2s_reg[21], pp_reg[116], r3c[19], r3s[20], r3c[20]);
FA	inst1108	(r2s_reg[22], pp_reg[117], r3c[20], r3s[21], r3c[21]);
FA	inst1109	(r2s_reg[23], pp_reg[118], r3c[21], r3s[22], r3c[22]);
FA	inst1110	(r2s_reg[24], pp_reg[119], r3c[22], r3s[23], r3c[23]);
FA	inst1111	(r2s_reg[25], pp_reg[120], r3c[23], r3s[24], r3c[24]);
FA	inst1112	(r2s_reg[26], pp_reg[121], r3c[24], r3s[25], r3c[25]);
FA	inst1113	(r2s_reg[27], pp_reg[122], r3c[25], r3s[26], r3c[26]);
FA	inst1114	(r2s_reg[28], pp_reg[123], r3c[26], r3s[27], r3c[27]);
FA	inst1115	(r2s_reg[29], pp_reg[124], r3c[27], r3s[28], r3c[28]);
FA	inst1116	(r2s_reg[30], pp_reg[94], r3c[28], r3s[29], r3c[29]);
FA	inst1117	(rc_last_reg[1], pp_reg[95], r3c[29], r3s[30], r3c[30]);
//Posible pipline
always @(posedge clk) begin
	r3s_reg <= r3s;
	rc_last_reg[2] <= r3c[30];
	ProcConditon_reg[3] <= ProcConditon_reg[2];
end

HA	inst1118	(r3s_reg[1], pp_reg[128], m[4], r4c[0]);
FA	inst1119	(r3s_reg[2], pp_reg[129], r4c[0], r4s[1], r4c[1]);
FA	inst1120	(r3s_reg[3], pp_reg[130], r4c[1], r4s[2], r4c[2]);
FA	inst1121	(r3s_reg[4], pp_reg[131], r4c[2], r4s[3], r4c[3]);
FA	inst1122	(r3s_reg[5], pp_reg[132], r4c[3], r4s[4], r4c[4]);
FA	inst1123	(r3s_reg[6], pp_reg[133], r4c[4], r4s[5], r4c[5]);
FA	inst1124	(r3s_reg[7], pp_reg[134], r4c[5], r4s[6], r4c[6]);
FA	inst1125	(r3s_reg[8], pp_reg[135], r4c[6], r4s[7], r4c[7]);
FA	inst1126	(r3s_reg[9], pp_reg[136], r4c[7], r4s[8], r4c[8]);
FA	inst1127	(r3s_reg[10], pp_reg[137], r4c[8], r4s[9], r4c[9]);
FA	inst1128	(r3s_reg[11], pp_reg[138], r4c[9], r4s[10], r4c[10]);
FA	inst1129	(r3s_reg[12], pp_reg[139], r4c[10], r4s[11], r4c[11]);
FA	inst1130	(r3s_reg[13], pp_reg[140], r4c[11], r4s[12], r4c[12]);
FA	inst1131	(r3s_reg[14], pp_reg[141], r4c[12], r4s[13], r4c[13]);
FA	inst1132	(r3s_reg[15], pp_reg[142], r4c[13], r4s[14], r4c[14]);
FA	inst1133	(r3s_reg[16], pp_reg[143], r4c[14], r4s[15], r4c[15]);
FA	inst1134	(r3s_reg[17], pp_reg[144], r4c[15], r4s[16], r4c[16]);
FA	inst1135	(r3s_reg[18], pp_reg[145], r4c[16], r4s[17], r4c[17]);
FA	inst1136	(r3s_reg[19], pp_reg[146], r4c[17], r4s[18], r4c[18]);
FA	inst1137	(r3s_reg[20], pp_reg[147], r4c[18], r4s[19], r4c[19]);
FA	inst1138	(r3s_reg[21], pp_reg[148], r4c[19], r4s[20], r4c[20]);
FA	inst1139	(r3s_reg[22], pp_reg[149], r4c[20], r4s[21], r4c[21]);
FA	inst1140	(r3s_reg[23], pp_reg[150], r4c[21], r4s[22], r4c[22]);
FA	inst1141	(r3s_reg[24], pp_reg[151], r4c[22], r4s[23], r4c[23]);
FA	inst1142	(r3s_reg[25], pp_reg[152], r4c[23], r4s[24], r4c[24]);
FA	inst1143	(r3s_reg[26], pp_reg[153], r4c[24], r4s[25], r4c[25]);
FA	inst1144	(r3s_reg[27], pp_reg[154], r4c[25], r4s[26], r4c[26]);
FA	inst1145	(r3s_reg[28], pp_reg[155], r4c[26], r4s[27], r4c[27]);
FA	inst1146	(r3s_reg[29], pp_reg[125], r4c[27], r4s[28], r4c[28]);
FA	inst1147	(r3s_reg[30], pp_reg[126], r4c[28], r4s[29], r4c[29]);
FA	inst1148	(rc_last_reg[2], pp_reg[127], r4c[29], r4s[30], r4c[30]);
//Posible pipline
always @(posedge clk) begin
	r4s_reg <= r4s;
	rc_last_reg[3] <= r4c[30];
	ProcConditon_reg[4] <= ProcConditon_reg[3];
end

HA	inst1149	(r4s_reg[1], pp_reg[160], m[5], r5c[0]);
FA	inst1150	(r4s_reg[2], pp_reg[161], r5c[0], r5s[1], r5c[1]);
FA	inst1151	(r4s_reg[3], pp_reg[162], r5c[1], r5s[2], r5c[2]);
FA	inst1152	(r4s_reg[4], pp_reg[163], r5c[2], r5s[3], r5c[3]);
FA	inst1153	(r4s_reg[5], pp_reg[164], r5c[3], r5s[4], r5c[4]);
FA	inst1154	(r4s_reg[6], pp_reg[165], r5c[4], r5s[5], r5c[5]);
FA	inst1155	(r4s_reg[7], pp_reg[166], r5c[5], r5s[6], r5c[6]);
FA	inst1156	(r4s_reg[8], pp_reg[167], r5c[6], r5s[7], r5c[7]);
FA	inst1157	(r4s_reg[9], pp_reg[168], r5c[7], r5s[8], r5c[8]);
FA	inst1158	(r4s_reg[10], pp_reg[169], r5c[8], r5s[9], r5c[9]);
FA	inst1159	(r4s_reg[11], pp_reg[170], r5c[9], r5s[10], r5c[10]);
FA	inst1160	(r4s_reg[12], pp_reg[171], r5c[10], r5s[11], r5c[11]);
FA	inst1161	(r4s_reg[13], pp_reg[172], r5c[11], r5s[12], r5c[12]);
FA	inst1162	(r4s_reg[14], pp_reg[173], r5c[12], r5s[13], r5c[13]);
FA	inst1163	(r4s_reg[15], pp_reg[174], r5c[13], r5s[14], r5c[14]);
FA	inst1164	(r4s_reg[16], pp_reg[175], r5c[14], r5s[15], r5c[15]);
FA	inst1165	(r4s_reg[17], pp_reg[176], r5c[15], r5s[16], r5c[16]);
FA	inst1166	(r4s_reg[18], pp_reg[177], r5c[16], r5s[17], r5c[17]);
FA	inst1167	(r4s_reg[19], pp_reg[178], r5c[17], r5s[18], r5c[18]);
FA	inst1168	(r4s_reg[20], pp_reg[179], r5c[18], r5s[19], r5c[19]);
FA	inst1169	(r4s_reg[21], pp_reg[180], r5c[19], r5s[20], r5c[20]);
FA	inst1170	(r4s_reg[22], pp_reg[181], r5c[20], r5s[21], r5c[21]);
FA	inst1171	(r4s_reg[23], pp_reg[182], r5c[21], r5s[22], r5c[22]);
FA	inst1172	(r4s_reg[24], pp_reg[183], r5c[22], r5s[23], r5c[23]);
FA	inst1173	(r4s_reg[25], pp_reg[184], r5c[23], r5s[24], r5c[24]);
FA	inst1174	(r4s_reg[26], pp_reg[185], r5c[24], r5s[25], r5c[25]);
FA	inst1175	(r4s_reg[27], pp_reg[186], r5c[25], r5s[26], r5c[26]);
FA	inst1176	(r4s_reg[28], pp_reg[156], r5c[26], r5s[27], r5c[27]);
FA	inst1177	(r4s_reg[29], pp_reg[157], r5c[27], r5s[28], r5c[28]);
FA	inst1178	(r4s_reg[30], pp_reg[158], r5c[28], r5s[29], r5c[29]);
FA	inst1179	(rc_last_reg[3], pp_reg[159], r5c[29], r5s[30], r5c[30]);
//Posible pipline

//Posible pipline
always @(posedge clk) begin
	r5s_reg <= r5s;
	rc_last_reg[4] <= r5c[30];
	ProcConditon_reg[5] <= ProcConditon_reg[4];
end

HA	inst1180	(r5s_reg[1], pp_reg[192], m[6], r6c[0]);
FA	inst1181	(r5s_reg[2], pp_reg[193], r6c[0], r6s[1], r6c[1]);
FA	inst1182	(r5s_reg[3], pp_reg[194], r6c[1], r6s[2], r6c[2]);
FA	inst1183	(r5s_reg[4], pp_reg[195], r6c[2], r6s[3], r6c[3]);
FA	inst1184	(r5s_reg[5], pp_reg[196], r6c[3], r6s[4], r6c[4]);
FA	inst1185	(r5s_reg[6], pp_reg[197], r6c[4], r6s[5], r6c[5]);
FA	inst1186	(r5s_reg[7], pp_reg[198], r6c[5], r6s[6], r6c[6]);
FA	inst1187	(r5s_reg[8], pp_reg[199], r6c[6], r6s[7], r6c[7]);
FA	inst1188	(r5s_reg[9], pp_reg[200], r6c[7], r6s[8], r6c[8]);
FA	inst1189	(r5s_reg[10], pp_reg[201], r6c[8], r6s[9], r6c[9]);
FA	inst1190	(r5s_reg[11], pp_reg[202], r6c[9], r6s[10], r6c[10]);
FA	inst1191	(r5s_reg[12], pp_reg[203], r6c[10], r6s[11], r6c[11]);
FA	inst1192	(r5s_reg[13], pp_reg[204], r6c[11], r6s[12], r6c[12]);
FA	inst1193	(r5s_reg[14], pp_reg[205], r6c[12], r6s[13], r6c[13]);
FA	inst1194	(r5s_reg[15], pp_reg[206], r6c[13], r6s[14], r6c[14]);
FA	inst1195	(r5s_reg[16], pp_reg[207], r6c[14], r6s[15], r6c[15]);
FA	inst1196	(r5s_reg[17], pp_reg[208], r6c[15], r6s[16], r6c[16]);
FA	inst1197	(r5s_reg[18], pp_reg[209], r6c[16], r6s[17], r6c[17]);
FA	inst1198	(r5s_reg[19], pp_reg[210], r6c[17], r6s[18], r6c[18]);
FA	inst1199	(r5s_reg[20], pp_reg[211], r6c[18], r6s[19], r6c[19]);
FA	inst1200	(r5s_reg[21], pp_reg[212], r6c[19], r6s[20], r6c[20]);
FA	inst1201	(r5s_reg[22], pp_reg[213], r6c[20], r6s[21], r6c[21]);
FA	inst1202	(r5s_reg[23], pp_reg[214], r6c[21], r6s[22], r6c[22]);
FA	inst1203	(r5s_reg[24], pp_reg[215], r6c[22], r6s[23], r6c[23]);
FA	inst1204	(r5s_reg[25], pp_reg[216], r6c[23], r6s[24], r6c[24]);
FA	inst1205	(r5s_reg[26], pp_reg[217], r6c[24], r6s[25], r6c[25]);
FA	inst1206	(r5s_reg[27], pp_reg[187], r6c[25], r6s[26], r6c[26]);
FA	inst1207	(r5s_reg[28], pp_reg[188], r6c[26], r6s[27], r6c[27]);
FA	inst1208	(r5s_reg[29], pp_reg[189], r6c[27], r6s[28], r6c[28]);
FA	inst1209	(r5s_reg[30], pp_reg[190], r6c[28], r6s[29], r6c[29]);
FA	inst1210	(rc_last_reg[4], pp_reg[191], r6c[29], r6s[30], r6c[30]);
//Posible pipline
always @(posedge clk) begin
	r6s_reg <= r6s;
	rc_last_reg[5] <= r6c[30];
	ProcConditon_reg[6] <= ProcConditon_reg[5];
end


HA	inst1211	(r6s_reg[1], pp_reg[224], m[7], r7c[0]);
FA	inst1212	(r6s_reg[2], pp_reg[225], r7c[0], r7s[1], r7c[1]);
FA	inst1213	(r6s_reg[3], pp_reg[226], r7c[1], r7s[2], r7c[2]);
FA	inst1214	(r6s_reg[4], pp_reg[227], r7c[2], r7s[3], r7c[3]);
FA	inst1215	(r6s_reg[5], pp_reg[228], r7c[3], r7s[4], r7c[4]);
FA	inst1216	(r6s_reg[6], pp_reg[229], r7c[4], r7s[5], r7c[5]);
FA	inst1217	(r6s_reg[7], pp_reg[230], r7c[5], r7s[6], r7c[6]);
FA	inst1218	(r6s_reg[8], pp_reg[231], r7c[6], r7s[7], r7c[7]);
FA	inst1219	(r6s_reg[9], pp_reg[232], r7c[7], r7s[8], r7c[8]);
FA	inst1220	(r6s_reg[10], pp_reg[233], r7c[8], r7s[9], r7c[9]);
FA	inst1221	(r6s_reg[11], pp_reg[234], r7c[9], r7s[10], r7c[10]);
FA	inst1222	(r6s_reg[12], pp_reg[235], r7c[10], r7s[11], r7c[11]);
FA	inst1223	(r6s_reg[13], pp_reg[236], r7c[11], r7s[12], r7c[12]);
FA	inst1224	(r6s_reg[14], pp_reg[237], r7c[12], r7s[13], r7c[13]);
FA	inst1225	(r6s_reg[15], pp_reg[238], r7c[13], r7s[14], r7c[14]);
FA	inst1226	(r6s_reg[16], pp_reg[239], r7c[14], r7s[15], r7c[15]);
FA	inst1227	(r6s_reg[17], pp_reg[240], r7c[15], r7s[16], r7c[16]);
FA	inst1228	(r6s_reg[18], pp_reg[241], r7c[16], r7s[17], r7c[17]);
FA	inst1229	(r6s_reg[19], pp_reg[242], r7c[17], r7s[18], r7c[18]);
FA	inst1230	(r6s_reg[20], pp_reg[243], r7c[18], r7s[19], r7c[19]);
FA	inst1231	(r6s_reg[21], pp_reg[244], r7c[19], r7s[20], r7c[20]);
FA	inst1232	(r6s_reg[22], pp_reg[245], r7c[20], r7s[21], r7c[21]);
FA	inst1233	(r6s_reg[23], pp_reg[246], r7c[21], r7s[22], r7c[22]);
FA	inst1234	(r6s_reg[24], pp_reg[247], r7c[22], r7s[23], r7c[23]);
FA	inst1235	(r6s_reg[25], pp_reg[248], r7c[23], r7s[24], r7c[24]);
FA	inst1236	(r6s_reg[26], pp_reg[218], r7c[24], r7s[25], r7c[25]);
FA	inst1237	(r6s_reg[27], pp_reg[219], r7c[25], r7s[26], r7c[26]);
FA	inst1238	(r6s_reg[28], pp_reg[220], r7c[26], r7s[27], r7c[27]);
FA	inst1239	(r6s_reg[29], pp_reg[221], r7c[27], r7s[28], r7c[28]);
FA	inst1240	(r6s_reg[30], pp_reg[222], r7c[28], r7s[29], r7c[29]);
FA	inst1241	(rc_last_reg[5], pp_reg[223], r7c[29], r7s[30], r7c[30]);
//Posible pipline
always @(posedge clk) begin
	r7s_reg <= r7s;
	rc_last_reg[6] <= r7c[30];
	ProcConditon_reg[7] <= ProcConditon_reg[6];
end

HA	inst1242	(r7s_reg[1], pp_reg[256], m[8], r8c[0]);
FA	inst1243	(r7s_reg[2], pp_reg[257], r8c[0], r8s[1], r8c[1]);
FA	inst1244	(r7s_reg[3], pp_reg[258], r8c[1], r8s[2], r8c[2]);
FA	inst1245	(r7s_reg[4], pp_reg[259], r8c[2], r8s[3], r8c[3]);
FA	inst1246	(r7s_reg[5], pp_reg[260], r8c[3], r8s[4], r8c[4]);
FA	inst1247	(r7s_reg[6], pp_reg[261], r8c[4], r8s[5], r8c[5]);
FA	inst1248	(r7s_reg[7], pp_reg[262], r8c[5], r8s[6], r8c[6]);
FA	inst1249	(r7s_reg[8], pp_reg[263], r8c[6], r8s[7], r8c[7]);
FA	inst1250	(r7s_reg[9], pp_reg[264], r8c[7], r8s[8], r8c[8]);
FA	inst1251	(r7s_reg[10], pp_reg[265], r8c[8], r8s[9], r8c[9]);
FA	inst1252	(r7s_reg[11], pp_reg[266], r8c[9], r8s[10], r8c[10]);
FA	inst1253	(r7s_reg[12], pp_reg[267], r8c[10], r8s[11], r8c[11]);
FA	inst1254	(r7s_reg[13], pp_reg[268], r8c[11], r8s[12], r8c[12]);
FA	inst1255	(r7s_reg[14], pp_reg[269], r8c[12], r8s[13], r8c[13]);
FA	inst1256	(r7s_reg[15], pp_reg[270], r8c[13], r8s[14], r8c[14]);
FA	inst1257	(r7s_reg[16], pp_reg[271], r8c[14], r8s[15], r8c[15]);
FA	inst1258	(r7s_reg[17], pp_reg[272], r8c[15], r8s[16], r8c[16]);
FA	inst1259	(r7s_reg[18], pp_reg[273], r8c[16], r8s[17], r8c[17]);
FA	inst1260	(r7s_reg[19], pp_reg[274], r8c[17], r8s[18], r8c[18]);
FA	inst1261	(r7s_reg[20], pp_reg[275], r8c[18], r8s[19], r8c[19]);
FA	inst1262	(r7s_reg[21], pp_reg[276], r8c[19], r8s[20], r8c[20]);
FA	inst1263	(r7s_reg[22], pp_reg[277], r8c[20], r8s[21], r8c[21]);
FA	inst1264	(r7s_reg[23], pp_reg[278], r8c[21], r8s[22], r8c[22]);
FA	inst1265	(r7s_reg[24], pp_reg[279], r8c[22], r8s[23], r8c[23]);
FA	inst1266	(r7s_reg[25], pp_reg[249], r8c[23], r8s[24], r8c[24]);
FA	inst1267	(r7s_reg[26], pp_reg[250], r8c[24], r8s[25], r8c[25]);
FA	inst1268	(r7s_reg[27], pp_reg[251], r8c[25], r8s[26], r8c[26]);
FA	inst1269	(r7s_reg[28], pp_reg[252], r8c[26], r8s[27], r8c[27]);
FA	inst1270	(r7s_reg[29], pp_reg[253], r8c[27], r8s[28], r8c[28]);
FA	inst1271	(r7s_reg[30], pp_reg[254], r8c[28], r8s[29], r8c[29]);
FA	inst1272	(rc_last_reg[6], pp_reg[255], r8c[29], r8s[30], r8c[30]);
//Posible pipline
always @(posedge clk) begin
	r8s_reg <= r8s;
	rc_last_reg[7] <= r8c[30];
	ProcConditon_reg[8] <= ProcConditon_reg[7];
end

HA	inst1273	(r8s_reg[1], pp_reg[288], m[9], r9c[0]);
FA	inst1274	(r8s_reg[2], pp_reg[289], r9c[0], r9s[1], r9c[1]);
FA	inst1275	(r8s_reg[3], pp_reg[290], r9c[1], r9s[2], r9c[2]);
FA	inst1276	(r8s_reg[4], pp_reg[291], r9c[2], r9s[3], r9c[3]);
FA	inst1277	(r8s_reg[5], pp_reg[292], r9c[3], r9s[4], r9c[4]);
FA	inst1278	(r8s_reg[6], pp_reg[293], r9c[4], r9s[5], r9c[5]);
FA	inst1279	(r8s_reg[7], pp_reg[294], r9c[5], r9s[6], r9c[6]);
FA	inst1280	(r8s_reg[8], pp_reg[295], r9c[6], r9s[7], r9c[7]);
FA	inst1281	(r8s_reg[9], pp_reg[296], r9c[7], r9s[8], r9c[8]);
FA	inst1282	(r8s_reg[10], pp_reg[297], r9c[8], r9s[9], r9c[9]);
FA	inst1283	(r8s_reg[11], pp_reg[298], r9c[9], r9s[10], r9c[10]);
FA	inst1284	(r8s_reg[12], pp_reg[299], r9c[10], r9s[11], r9c[11]);
FA	inst1285	(r8s_reg[13], pp_reg[300], r9c[11], r9s[12], r9c[12]);
FA	inst1286	(r8s_reg[14], pp_reg[301], r9c[12], r9s[13], r9c[13]);
FA	inst1287	(r8s_reg[15], pp_reg[302], r9c[13], r9s[14], r9c[14]);
FA	inst1288	(r8s_reg[16], pp_reg[303], r9c[14], r9s[15], r9c[15]);
FA	inst1289	(r8s_reg[17], pp_reg[304], r9c[15], r9s[16], r9c[16]);
FA	inst1290	(r8s_reg[18], pp_reg[305], r9c[16], r9s[17], r9c[17]);
FA	inst1291	(r8s_reg[19], pp_reg[306], r9c[17], r9s[18], r9c[18]);
FA	inst1292	(r8s_reg[20], pp_reg[307], r9c[18], r9s[19], r9c[19]);
FA	inst1293	(r8s_reg[21], pp_reg[308], r9c[19], r9s[20], r9c[20]);
FA	inst1294	(r8s_reg[22], pp_reg[309], r9c[20], r9s[21], r9c[21]);
FA	inst1295	(r8s_reg[23], pp_reg[310], r9c[21], r9s[22], r9c[22]);
FA	inst1296	(r8s_reg[24], pp_reg[280], r9c[22], r9s[23], r9c[23]);
FA	inst1297	(r8s_reg[25], pp_reg[281], r9c[23], r9s[24], r9c[24]);
FA	inst1298	(r8s_reg[26], pp_reg[282], r9c[24], r9s[25], r9c[25]);
FA	inst1299	(r8s_reg[27], pp_reg[283], r9c[25], r9s[26], r9c[26]);
FA	inst1300	(r8s_reg[28], pp_reg[284], r9c[26], r9s[27], r9c[27]);
FA	inst1301	(r8s_reg[29], pp_reg[285], r9c[27], r9s[28], r9c[28]);
FA	inst1302	(r8s_reg[30], pp_reg[286], r9c[28], r9s[29], r9c[29]);
FA	inst1303	(rc_last_reg[7], pp_reg[287], r9c[29], r9s[30], r9c[30]);
//Posible pipline

always @(posedge clk) begin
	r9s_reg <= r9s;
	rc_last_reg[8] <= r9c[30];
	ProcConditon_reg[9] <= ProcConditon_reg[8];
end

HA	inst1304	(r9s_reg[1], pp_reg[320], m[10], r10c[0]);
FA	inst1305	(r9s_reg[2], pp_reg[321], r10c[0], r10s[1], r10c[1]);
FA	inst1306	(r9s_reg[3], pp_reg[322], r10c[1], r10s[2], r10c[2]);
FA	inst1307	(r9s_reg[4], pp_reg[323], r10c[2], r10s[3], r10c[3]);
FA	inst1308	(r9s_reg[5], pp_reg[324], r10c[3], r10s[4], r10c[4]);
FA	inst1309	(r9s_reg[6], pp_reg[325], r10c[4], r10s[5], r10c[5]);
FA	inst1310	(r9s_reg[7], pp_reg[326], r10c[5], r10s[6], r10c[6]);
FA	inst1311	(r9s_reg[8], pp_reg[327], r10c[6], r10s[7], r10c[7]);
FA	inst1312	(r9s_reg[9], pp_reg[328], r10c[7], r10s[8], r10c[8]);
FA	inst1313	(r9s_reg[10], pp_reg[329], r10c[8], r10s[9], r10c[9]);
FA	inst1314	(r9s_reg[11], pp_reg[330], r10c[9], r10s[10], r10c[10]);
FA	inst1315	(r9s_reg[12], pp_reg[331], r10c[10], r10s[11], r10c[11]);
FA	inst1316	(r9s_reg[13], pp_reg[332], r10c[11], r10s[12], r10c[12]);
FA	inst1317	(r9s_reg[14], pp_reg[333], r10c[12], r10s[13], r10c[13]);
FA	inst1318	(r9s_reg[15], pp_reg[334], r10c[13], r10s[14], r10c[14]);
FA	inst1319	(r9s_reg[16], pp_reg[335], r10c[14], r10s[15], r10c[15]);
FA	inst1320	(r9s_reg[17], pp_reg[336], r10c[15], r10s[16], r10c[16]);
FA	inst1321	(r9s_reg[18], pp_reg[337], r10c[16], r10s[17], r10c[17]);
FA	inst1322	(r9s_reg[19], pp_reg[338], r10c[17], r10s[18], r10c[18]);
FA	inst1323	(r9s_reg[20], pp_reg[339], r10c[18], r10s[19], r10c[19]);
FA	inst1324	(r9s_reg[21], pp_reg[340], r10c[19], r10s[20], r10c[20]);
FA	inst1325	(r9s_reg[22], pp_reg[341], r10c[20], r10s[21], r10c[21]);
FA	inst1326	(r9s_reg[23], pp_reg[311], r10c[21], r10s[22], r10c[22]);
FA	inst1327	(r9s_reg[24], pp_reg[312], r10c[22], r10s[23], r10c[23]);
FA	inst1328	(r9s_reg[25], pp_reg[313], r10c[23], r10s[24], r10c[24]);
FA	inst1329	(r9s_reg[26], pp_reg[314], r10c[24], r10s[25], r10c[25]);
FA	inst1330	(r9s_reg[27], pp_reg[315], r10c[25], r10s[26], r10c[26]);
FA	inst1331	(r9s_reg[28], pp_reg[316], r10c[26], r10s[27], r10c[27]);
FA	inst1332	(r9s_reg[29], pp_reg[317], r10c[27], r10s[28], r10c[28]);
FA	inst1333	(r9s_reg[30], pp_reg[318], r10c[28], r10s[29], r10c[29]);
FA	inst1334	(rc_last_reg[8], pp_reg[319], r10c[29], r10s[30], r10c[30]);
//Posible pipline

always @(posedge clk) begin
	r10s_reg <= r10s;
	rc_last_reg[9] <= r10c[30];
	ProcConditon_reg[10] <= ProcConditon_reg[9];
end

HA	inst1335	(r10s_reg[1], pp_reg[352], m[11], r11c[0]);
FA	inst1336	(r10s_reg[2], pp_reg[353], r11c[0], r11s[1], r11c[1]);
FA	inst1337	(r10s_reg[3], pp_reg[354], r11c[1], r11s[2], r11c[2]);
FA	inst1338	(r10s_reg[4], pp_reg[355], r11c[2], r11s[3], r11c[3]);
FA	inst1339	(r10s_reg[5], pp_reg[356], r11c[3], r11s[4], r11c[4]);
FA	inst1340	(r10s_reg[6], pp_reg[357], r11c[4], r11s[5], r11c[5]);
FA	inst1341	(r10s_reg[7], pp_reg[358], r11c[5], r11s[6], r11c[6]);
FA	inst1342	(r10s_reg[8], pp_reg[359], r11c[6], r11s[7], r11c[7]);
FA	inst1343	(r10s_reg[9], pp_reg[360], r11c[7], r11s[8], r11c[8]);
FA	inst1344	(r10s_reg[10], pp_reg[361], r11c[8], r11s[9], r11c[9]);
FA	inst1345	(r10s_reg[11], pp_reg[362], r11c[9], r11s[10], r11c[10]);
FA	inst1346	(r10s_reg[12], pp_reg[363], r11c[10], r11s[11], r11c[11]);
FA	inst1347	(r10s_reg[13], pp_reg[364], r11c[11], r11s[12], r11c[12]);
FA	inst1348	(r10s_reg[14], pp_reg[365], r11c[12], r11s[13], r11c[13]);
FA	inst1349	(r10s_reg[15], pp_reg[366], r11c[13], r11s[14], r11c[14]);
FA	inst1350	(r10s_reg[16], pp_reg[367], r11c[14], r11s[15], r11c[15]);
FA	inst1351	(r10s_reg[17], pp_reg[368], r11c[15], r11s[16], r11c[16]);
FA	inst1352	(r10s_reg[18], pp_reg[369], r11c[16], r11s[17], r11c[17]);
FA	inst1353	(r10s_reg[19], pp_reg[370], r11c[17], r11s[18], r11c[18]);
FA	inst1354	(r10s_reg[20], pp_reg[371], r11c[18], r11s[19], r11c[19]);
FA	inst1355	(r10s_reg[21], pp_reg[372], r11c[19], r11s[20], r11c[20]);
FA	inst1356	(r10s_reg[22], pp_reg[342], r11c[20], r11s[21], r11c[21]);
FA	inst1357	(r10s_reg[23], pp_reg[343], r11c[21], r11s[22], r11c[22]);
FA	inst1358	(r10s_reg[24], pp_reg[344], r11c[22], r11s[23], r11c[23]);
FA	inst1359	(r10s_reg[25], pp_reg[345], r11c[23], r11s[24], r11c[24]);
FA	inst1360	(r10s_reg[26], pp_reg[346], r11c[24], r11s[25], r11c[25]);
FA	inst1361	(r10s_reg[27], pp_reg[347], r11c[25], r11s[26], r11c[26]);
FA	inst1362	(r10s_reg[28], pp_reg[348], r11c[26], r11s[27], r11c[27]);
FA	inst1363	(r10s_reg[29], pp_reg[349], r11c[27], r11s[28], r11c[28]);
FA	inst1364	(r10s_reg[30], pp_reg[350], r11c[28], r11s[29], r11c[29]);
FA	inst1365	(rc_last_reg[9], pp_reg[351], r11c[29], r11s[30], r11c[30]);
//Posible pipline
always @(posedge clk) begin
	r11s_reg <= r11s;
	rc_last_reg[10] <= r11c[30];
	ProcConditon_reg[11] <= ProcConditon_reg[10];
end

HA	inst1366	(r11s_reg[1], pp_reg[384], m[12], r12c[0]);
FA	inst1367	(r11s_reg[2], pp_reg[385], r12c[0], r12s[1], r12c[1]);
FA	inst1368	(r11s_reg[3], pp_reg[386], r12c[1], r12s[2], r12c[2]);
FA	inst1369	(r11s_reg[4], pp_reg[387], r12c[2], r12s[3], r12c[3]);
FA	inst1370	(r11s_reg[5], pp_reg[388], r12c[3], r12s[4], r12c[4]);
FA	inst1371	(r11s_reg[6], pp_reg[389], r12c[4], r12s[5], r12c[5]);
FA	inst1372	(r11s_reg[7], pp_reg[390], r12c[5], r12s[6], r12c[6]);
FA	inst1373	(r11s_reg[8], pp_reg[391], r12c[6], r12s[7], r12c[7]);
FA	inst1374	(r11s_reg[9], pp_reg[392], r12c[7], r12s[8], r12c[8]);
FA	inst1375	(r11s_reg[10], pp_reg[393], r12c[8], r12s[9], r12c[9]);
FA	inst1376	(r11s_reg[11], pp_reg[394], r12c[9], r12s[10], r12c[10]);
FA	inst1377	(r11s_reg[12], pp_reg[395], r12c[10], r12s[11], r12c[11]);
FA	inst1378	(r11s_reg[13], pp_reg[396], r12c[11], r12s[12], r12c[12]);
FA	inst1379	(r11s_reg[14], pp_reg[397], r12c[12], r12s[13], r12c[13]);
FA	inst1380	(r11s_reg[15], pp_reg[398], r12c[13], r12s[14], r12c[14]);
FA	inst1381	(r11s_reg[16], pp_reg[399], r12c[14], r12s[15], r12c[15]);
FA	inst1382	(r11s_reg[17], pp_reg[400], r12c[15], r12s[16], r12c[16]);
FA	inst1383	(r11s_reg[18], pp_reg[401], r12c[16], r12s[17], r12c[17]);
FA	inst1384	(r11s_reg[19], pp_reg[402], r12c[17], r12s[18], r12c[18]);
FA	inst1385	(r11s_reg[20], pp_reg[403], r12c[18], r12s[19], r12c[19]);
FA	inst1386	(r11s_reg[21], pp_reg[373], r12c[19], r12s[20], r12c[20]);
FA	inst1387	(r11s_reg[22], pp_reg[374], r12c[20], r12s[21], r12c[21]);
FA	inst1388	(r11s_reg[23], pp_reg[375], r12c[21], r12s[22], r12c[22]);
FA	inst1389	(r11s_reg[24], pp_reg[376], r12c[22], r12s[23], r12c[23]);
FA	inst1390	(r11s_reg[25], pp_reg[377], r12c[23], r12s[24], r12c[24]);
FA	inst1391	(r11s_reg[26], pp_reg[378], r12c[24], r12s[25], r12c[25]);
FA	inst1392	(r11s_reg[27], pp_reg[379], r12c[25], r12s[26], r12c[26]);
FA	inst1393	(r11s_reg[28], pp_reg[380], r12c[26], r12s[27], r12c[27]);
FA	inst1394	(r11s_reg[29], pp_reg[381], r12c[27], r12s[28], r12c[28]);
FA	inst1395	(r11s_reg[30], pp_reg[382], r12c[28], r12s[29], r12c[29]);
FA	inst1396	(rc_last_reg[10], pp_reg[383], r12c[29], r12s[30], r12c[30]);
//Posible pipline
always @(posedge clk) begin
	r12s_reg <= r12s;
	rc_last_reg[11] <= r12c[30];
	ProcConditon_reg[12] <= ProcConditon_reg[11];
end

HA	inst1397	(r12s_reg[1], pp_reg[416], m[13], r13c[0]);
FA	inst1398	(r12s_reg[2], pp_reg[417], r13c[0], r13s[1], r13c[1]);
FA	inst1399	(r12s_reg[3], pp_reg[418], r13c[1], r13s[2], r13c[2]);
FA	inst1400	(r12s_reg[4], pp_reg[419], r13c[2], r13s[3], r13c[3]);
FA	inst1401	(r12s_reg[5], pp_reg[420], r13c[3], r13s[4], r13c[4]);
FA	inst1402	(r12s_reg[6], pp_reg[421], r13c[4], r13s[5], r13c[5]);
FA	inst1403	(r12s_reg[7], pp_reg[422], r13c[5], r13s[6], r13c[6]);
FA	inst1404	(r12s_reg[8], pp_reg[423], r13c[6], r13s[7], r13c[7]);
FA	inst1405	(r12s_reg[9], pp_reg[424], r13c[7], r13s[8], r13c[8]);
FA	inst1406	(r12s_reg[10], pp_reg[425], r13c[8], r13s[9], r13c[9]);
FA	inst1407	(r12s_reg[11], pp_reg[426], r13c[9], r13s[10], r13c[10]);
FA	inst1408	(r12s_reg[12], pp_reg[427], r13c[10], r13s[11], r13c[11]);
FA	inst1409	(r12s_reg[13], pp_reg[428], r13c[11], r13s[12], r13c[12]);
FA	inst1410	(r12s_reg[14], pp_reg[429], r13c[12], r13s[13], r13c[13]);
FA	inst1411	(r12s_reg[15], pp_reg[430], r13c[13], r13s[14], r13c[14]);
FA	inst1412	(r12s_reg[16], pp_reg[431], r13c[14], r13s[15], r13c[15]);
FA	inst1413	(r12s_reg[17], pp_reg[432], r13c[15], r13s[16], r13c[16]);
FA	inst1414	(r12s_reg[18], pp_reg[433], r13c[16], r13s[17], r13c[17]);
FA	inst1415	(r12s_reg[19], pp_reg[434], r13c[17], r13s[18], r13c[18]);
FA	inst1416	(r12s_reg[20], pp_reg[404], r13c[18], r13s[19], r13c[19]);
FA	inst1417	(r12s_reg[21], pp_reg[405], r13c[19], r13s[20], r13c[20]);
FA	inst1418	(r12s_reg[22], pp_reg[406], r13c[20], r13s[21], r13c[21]);
FA	inst1419	(r12s_reg[23], pp_reg[407], r13c[21], r13s[22], r13c[22]);
FA	inst1420	(r12s_reg[24], pp_reg[408], r13c[22], r13s[23], r13c[23]);
FA	inst1421	(r12s_reg[25], pp_reg[409], r13c[23], r13s[24], r13c[24]);
FA	inst1422	(r12s_reg[26], pp_reg[410], r13c[24], r13s[25], r13c[25]);
FA	inst1423	(r12s_reg[27], pp_reg[411], r13c[25], r13s[26], r13c[26]);
FA	inst1424	(r12s_reg[28], pp_reg[412], r13c[26], r13s[27], r13c[27]);
FA	inst1425	(r12s_reg[29], pp_reg[413], r13c[27], r13s[28], r13c[28]);
FA	inst1426	(r12s_reg[30], pp_reg[414], r13c[28], r13s[29], r13c[29]);
FA	inst1427	(rc_last_reg[11], pp_reg[415], r13c[29], r13s[30], r13c[30]);
//Posible pipline
always @(posedge clk) begin
	r13s_reg <= r13s;
	rc_last_reg[12] <= r13c[30];
	ProcConditon_reg[13] <= ProcConditon_reg[12];
end


HA	inst1428	(r13s_reg[1], pp_reg[448], m[14], r14c[0]);
FA	inst1429	(r13s_reg[2], pp_reg[449], r14c[0], r14s[1], r14c[1]);
FA	inst1430	(r13s_reg[3], pp_reg[450], r14c[1], r14s[2], r14c[2]);
FA	inst1431	(r13s_reg[4], pp_reg[451], r14c[2], r14s[3], r14c[3]);
FA	inst1432	(r13s_reg[5], pp_reg[452], r14c[3], r14s[4], r14c[4]);
FA	inst1433	(r13s_reg[6], pp_reg[453], r14c[4], r14s[5], r14c[5]);
FA	inst1434	(r13s_reg[7], pp_reg[454], r14c[5], r14s[6], r14c[6]);
FA	inst1435	(r13s_reg[8], pp_reg[455], r14c[6], r14s[7], r14c[7]);
FA	inst1436	(r13s_reg[9], pp_reg[456], r14c[7], r14s[8], r14c[8]);
FA	inst1437	(r13s_reg[10], pp_reg[457], r14c[8], r14s[9], r14c[9]);
FA	inst1438	(r13s_reg[11], pp_reg[458], r14c[9], r14s[10], r14c[10]);
FA	inst1439	(r13s_reg[12], pp_reg[459], r14c[10], r14s[11], r14c[11]);
FA	inst1440	(r13s_reg[13], pp_reg[460], r14c[11], r14s[12], r14c[12]);
FA	inst1441	(r13s_reg[14], pp_reg[461], r14c[12], r14s[13], r14c[13]);
FA	inst1442	(r13s_reg[15], pp_reg[462], r14c[13], r14s[14], r14c[14]);
FA	inst1443	(r13s_reg[16], pp_reg[463], r14c[14], r14s[15], r14c[15]);
FA	inst1444	(r13s_reg[17], pp_reg[464], r14c[15], r14s[16], r14c[16]);
FA	inst1445	(r13s_reg[18], pp_reg[465], r14c[16], r14s[17], r14c[17]);
FA	inst1446	(r13s_reg[19], pp_reg[435], r14c[17], r14s[18], r14c[18]);
FA	inst1447	(r13s_reg[20], pp_reg[436], r14c[18], r14s[19], r14c[19]);
FA	inst1448	(r13s_reg[21], pp_reg[437], r14c[19], r14s[20], r14c[20]);
FA	inst1449	(r13s_reg[22], pp_reg[438], r14c[20], r14s[21], r14c[21]);
FA	inst1450	(r13s_reg[23], pp_reg[439], r14c[21], r14s[22], r14c[22]);
FA	inst1451	(r13s_reg[24], pp_reg[440], r14c[22], r14s[23], r14c[23]);
FA	inst1452	(r13s_reg[25], pp_reg[441], r14c[23], r14s[24], r14c[24]);
FA	inst1453	(r13s_reg[26], pp_reg[442], r14c[24], r14s[25], r14c[25]);
FA	inst1454	(r13s_reg[27], pp_reg[443], r14c[25], r14s[26], r14c[26]);
FA	inst1455	(r13s_reg[28], pp_reg[444], r14c[26], r14s[27], r14c[27]);
FA	inst1456	(r13s_reg[29], pp_reg[445], r14c[27], r14s[28], r14c[28]);
FA	inst1457	(r13s_reg[30], pp_reg[446], r14c[28], r14s[29], r14c[29]);
FA	inst1458	(rc_last_reg[12], pp_reg[447], r14c[29], r14s[30], r14c[30]);
//Posible pipline
always @(posedge clk) begin
	r14s_reg <= r14s;
	rc_last_reg[13] <= r14c[30];
	ProcConditon_reg[14] <= ProcConditon_reg[13];
end



HA	inst1459	(r14s_reg[1], pp_reg[480], m[15], r15c[0]);
FA	inst1460	(r14s_reg[2], pp_reg[481], r15c[0], r15s[1], r15c[1]);
FA	inst1461	(r14s_reg[3], pp_reg[482], r15c[1], r15s[2], r15c[2]);
FA	inst1462	(r14s_reg[4], pp_reg[483], r15c[2], r15s[3], r15c[3]);
FA	inst1463	(r14s_reg[5], pp_reg[484], r15c[3], r15s[4], r15c[4]);
FA	inst1464	(r14s_reg[6], pp_reg[485], r15c[4], r15s[5], r15c[5]);
FA	inst1465	(r14s_reg[7], pp_reg[486], r15c[5], r15s[6], r15c[6]);
FA	inst1466	(r14s_reg[8], pp_reg[487], r15c[6], r15s[7], r15c[7]);
FA	inst1467	(r14s_reg[9], pp_reg[488], r15c[7], r15s[8], r15c[8]);
FA	inst1468	(r14s_reg[10], pp_reg[489], r15c[8], r15s[9], r15c[9]);
FA	inst1469	(r14s_reg[11], pp_reg[490], r15c[9], r15s[10], r15c[10]);
FA	inst1470	(r14s_reg[12], pp_reg[491], r15c[10], r15s[11], r15c[11]);
FA	inst1471	(r14s_reg[13], pp_reg[492], r15c[11], r15s[12], r15c[12]);
FA	inst1472	(r14s_reg[14], pp_reg[493], r15c[12], r15s[13], r15c[13]);
FA	inst1473	(r14s_reg[15], pp_reg[494], r15c[13], r15s[14], r15c[14]);
FA	inst1474	(r14s_reg[16], pp_reg[495], r15c[14], r15s[15], r15c[15]);
FA	inst1475	(r14s_reg[17], pp_reg[496], r15c[15], r15s[16], r15c[16]);
FA	inst1476	(r14s_reg[18], pp_reg[466], r15c[16], r15s[17], r15c[17]);
FA	inst1477	(r14s_reg[19], pp_reg[467], r15c[17], r15s[18], r15c[18]);
FA	inst1478	(r14s_reg[20], pp_reg[468], r15c[18], r15s[19], r15c[19]);
FA	inst1479	(r14s_reg[21], pp_reg[469], r15c[19], r15s[20], r15c[20]);
FA	inst1480	(r14s_reg[22], pp_reg[470], r15c[20], r15s[21], r15c[21]);
FA	inst1481	(r14s_reg[23], pp_reg[471], r15c[21], r15s[22], r15c[22]);
FA	inst1482	(r14s_reg[24], pp_reg[472], r15c[22], r15s[23], r15c[23]);
FA	inst1483	(r14s_reg[25], pp_reg[473], r15c[23], r15s[24], r15c[24]);
FA	inst1484	(r14s_reg[26], pp_reg[474], r15c[24], r15s[25], r15c[25]);
FA	inst1485	(r14s_reg[27], pp_reg[475], r15c[25], r15s[26], r15c[26]);
FA	inst1486	(r14s_reg[28], pp_reg[476], r15c[26], r15s[27], r15c[27]);
FA	inst1487	(r14s_reg[29], pp_reg[477], r15c[27], r15s[28], r15c[28]);
FA	inst1488	(r14s_reg[30], pp_reg[478], r15c[28], r15s[29], r15c[29]);
FA	inst1489	(rc_last_reg[13], pp_reg[479], r15c[29], r15s[30], r15c[30]);
//Posible pipline
always @(posedge clk) begin
	r15s_reg <= r15s;
	rc_last_reg[14] <= r15c[30];
	ProcConditon_reg[15] <= ProcConditon_reg[14];
end

HA	inst1490	(r15s_reg[1], pp_reg[512], m[16], r16c[0]);
FA	inst1491	(r15s_reg[2], pp_reg[513], r16c[0], r16s[1], r16c[1]);
FA	inst1492	(r15s_reg[3], pp_reg[514], r16c[1], r16s[2], r16c[2]);
FA	inst1493	(r15s_reg[4], pp_reg[515], r16c[2], r16s[3], r16c[3]);
FA	inst1494	(r15s_reg[5], pp_reg[516], r16c[3], r16s[4], r16c[4]);
FA	inst1495	(r15s_reg[6], pp_reg[517], r16c[4], r16s[5], r16c[5]);
FA	inst1496	(r15s_reg[7], pp_reg[518], r16c[5], r16s[6], r16c[6]);
FA	inst1497	(r15s_reg[8], pp_reg[519], r16c[6], r16s[7], r16c[7]);
FA	inst1498	(r15s_reg[9], pp_reg[520], r16c[7], r16s[8], r16c[8]);
FA	inst1499	(r15s_reg[10], pp_reg[521], r16c[8], r16s[9], r16c[9]);
FA	inst1500	(r15s_reg[11], pp_reg[522], r16c[9], r16s[10], r16c[10]);
FA	inst1501	(r15s_reg[12], pp_reg[523], r16c[10], r16s[11], r16c[11]);
FA	inst1502	(r15s_reg[13], pp_reg[524], r16c[11], r16s[12], r16c[12]);
FA	inst1503	(r15s_reg[14], pp_reg[525], r16c[12], r16s[13], r16c[13]);
FA	inst1504	(r15s_reg[15], pp_reg[526], r16c[13], r16s[14], r16c[14]);
FA	inst1505	(r15s_reg[16], pp_reg[527], r16c[14], r16s[15], r16c[15]);
FA	inst1506	(r15s_reg[17], pp_reg[497], r16c[15], r16s[16], r16c[16]);
FA	inst1507	(r15s_reg[18], pp_reg[498], r16c[16], r16s[17], r16c[17]);
FA	inst1508	(r15s_reg[19], pp_reg[499], r16c[17], r16s[18], r16c[18]);
FA	inst1509	(r15s_reg[20], pp_reg[500], r16c[18], r16s[19], r16c[19]);
FA	inst1510	(r15s_reg[21], pp_reg[501], r16c[19], r16s[20], r16c[20]);
FA	inst1511	(r15s_reg[22], pp_reg[502], r16c[20], r16s[21], r16c[21]);
FA	inst1512	(r15s_reg[23], pp_reg[503], r16c[21], r16s[22], r16c[22]);
FA	inst1513	(r15s_reg[24], pp_reg[504], r16c[22], r16s[23], r16c[23]);
FA	inst1514	(r15s_reg[25], pp_reg[505], r16c[23], r16s[24], r16c[24]);
FA	inst1515	(r15s_reg[26], pp_reg[506], r16c[24], r16s[25], r16c[25]);
FA	inst1516	(r15s_reg[27], pp_reg[507], r16c[25], r16s[26], r16c[26]);
FA	inst1517	(r15s_reg[28], pp_reg[508], r16c[26], r16s[27], r16c[27]);
FA	inst1518	(r15s_reg[29], pp_reg[509], r16c[27], r16s[28], r16c[28]);
FA	inst1519	(r15s_reg[30], pp_reg[510], r16c[28], r16s[29], r16c[29]);
FA	inst1520	(rc_last_reg[10], pp_reg[511], r16c[29], r16s[30], r16c[30]);
//Posible pipline
always @(posedge clk) begin
	r16s_reg <= r16s;
	rc_last_reg[15] <= r16c[30];
	ProcConditon_reg[16] <= ProcConditon_reg[15];
end

HA	inst1521	(r16s_reg[1], pp_reg[544], m[17], r17c[0]);
FA	inst1522	(r16s_reg[2], pp_reg[545], r17c[0], r17s[1], r17c[1]);
FA	inst1523	(r16s_reg[3], pp_reg[546], r17c[1], r17s[2], r17c[2]);
FA	inst1524	(r16s_reg[4], pp_reg[547], r17c[2], r17s[3], r17c[3]);
FA	inst1525	(r16s_reg[5], pp_reg[548], r17c[3], r17s[4], r17c[4]);
FA	inst1526	(r16s_reg[6], pp_reg[549], r17c[4], r17s[5], r17c[5]);
FA	inst1527	(r16s_reg[7], pp_reg[550], r17c[5], r17s[6], r17c[6]);
FA	inst1528	(r16s_reg[8], pp_reg[551], r17c[6], r17s[7], r17c[7]);
FA	inst1529	(r16s_reg[9], pp_reg[552], r17c[7], r17s[8], r17c[8]);
FA	inst1530	(r16s_reg[10], pp_reg[553], r17c[8], r17s[9], r17c[9]);
FA	inst1531	(r16s_reg[11], pp_reg[554], r17c[9], r17s[10], r17c[10]);
FA	inst1532	(r16s_reg[12], pp_reg[555], r17c[10], r17s[11], r17c[11]);
FA	inst1533	(r16s_reg[13], pp_reg[556], r17c[11], r17s[12], r17c[12]);
FA	inst1534	(r16s_reg[14], pp_reg[557], r17c[12], r17s[13], r17c[13]);
FA	inst1535	(r16s_reg[15], pp_reg[558], r17c[13], r17s[14], r17c[14]);
FA	inst1536	(r16s_reg[16], pp_reg[528], r17c[14], r17s[15], r17c[15]);
FA	inst1537	(r16s_reg[17], pp_reg[529], r17c[15], r17s[16], r17c[16]);
FA	inst1538	(r16s_reg[18], pp_reg[530], r17c[16], r17s[17], r17c[17]);
FA	inst1539	(r16s_reg[19], pp_reg[531], r17c[17], r17s[18], r17c[18]);
FA	inst1540	(r16s_reg[20], pp_reg[532], r17c[18], r17s[19], r17c[19]);
FA	inst1541	(r16s_reg[21], pp_reg[533], r17c[19], r17s[20], r17c[20]);
FA	inst1542	(r16s_reg[22], pp_reg[534], r17c[20], r17s[21], r17c[21]);
FA	inst1543	(r16s_reg[23], pp_reg[535], r17c[21], r17s[22], r17c[22]);
FA	inst1544	(r16s_reg[24], pp_reg[536], r17c[22], r17s[23], r17c[23]);
FA	inst1545	(r16s_reg[25], pp_reg[537], r17c[23], r17s[24], r17c[24]);
FA	inst1546	(r16s_reg[26], pp_reg[538], r17c[24], r17s[25], r17c[25]);
FA	inst1547	(r16s_reg[27], pp_reg[539], r17c[25], r17s[26], r17c[26]);
FA	inst1548	(r16s_reg[28], pp_reg[540], r17c[26], r17s[27], r17c[27]);
FA	inst1549	(r16s_reg[29], pp_reg[541], r17c[27], r17s[28], r17c[28]);
FA	inst1550	(r16s_reg[30], pp_reg[542], r17c[28], r17s[29], r17c[29]);
FA	inst1551	(rc_last_reg[15], pp_reg[543], r17c[29], r17s[30], r17c[30]);
//Posible pipline
always @(posedge clk) begin
	r17s_reg <= r17s;
	rc_last_reg[16] <= r17c[30];
	ProcConditon_reg[17] <= ProcConditon_reg[16];
end

HA	inst1552	(r17s_reg[1], pp_reg[576], m[18], r18c[0]);
FA	inst1553	(r17s_reg[2], pp_reg[577], r18c[0], r18s[1], r18c[1]);
FA	inst1554	(r17s_reg[3], pp_reg[578], r18c[1], r18s[2], r18c[2]);
FA	inst1555	(r17s_reg[4], pp_reg[579], r18c[2], r18s[3], r18c[3]);
FA	inst1556	(r17s_reg[5], pp_reg[580], r18c[3], r18s[4], r18c[4]);
FA	inst1557	(r17s_reg[6], pp_reg[581], r18c[4], r18s[5], r18c[5]);
FA	inst1558	(r17s_reg[7], pp_reg[582], r18c[5], r18s[6], r18c[6]);
FA	inst1559	(r17s_reg[8], pp_reg[583], r18c[6], r18s[7], r18c[7]);
FA	inst1560	(r17s_reg[9], pp_reg[584], r18c[7], r18s[8], r18c[8]);
FA	inst1561	(r17s_reg[10], pp_reg[585], r18c[8], r18s[9], r18c[9]);
FA	inst1562	(r17s_reg[11], pp_reg[586], r18c[9], r18s[10], r18c[10]);
FA	inst1563	(r17s_reg[12], pp_reg[587], r18c[10], r18s[11], r18c[11]);
FA	inst1564	(r17s_reg[13], pp_reg[588], r18c[11], r18s[12], r18c[12]);
FA	inst1565	(r17s_reg[14], pp_reg[589], r18c[12], r18s[13], r18c[13]);
FA	inst1566	(r17s_reg[15], pp_reg[559], r18c[13], r18s[14], r18c[14]);
FA	inst1567	(r17s_reg[16], pp_reg[560], r18c[14], r18s[15], r18c[15]);
FA	inst1568	(r17s_reg[17], pp_reg[561], r18c[15], r18s[16], r18c[16]);
FA	inst1569	(r17s_reg[18], pp_reg[562], r18c[16], r18s[17], r18c[17]);
FA	inst1570	(r17s_reg[19], pp_reg[563], r18c[17], r18s[18], r18c[18]);
FA	inst1571	(r17s_reg[20], pp_reg[564], r18c[18], r18s[19], r18c[19]);
FA	inst1572	(r17s_reg[21], pp_reg[565], r18c[19], r18s[20], r18c[20]);
FA	inst1573	(r17s_reg[22], pp_reg[566], r18c[20], r18s[21], r18c[21]);
FA	inst1574	(r17s_reg[23], pp_reg[567], r18c[21], r18s[22], r18c[22]);
FA	inst1575	(r17s_reg[24], pp_reg[568], r18c[22], r18s[23], r18c[23]);
FA	inst1576	(r17s_reg[25], pp_reg[569], r18c[23], r18s[24], r18c[24]);
FA	inst1577	(r17s_reg[26], pp_reg[570], r18c[24], r18s[25], r18c[25]);
FA	inst1578	(r17s_reg[27], pp_reg[571], r18c[25], r18s[26], r18c[26]);
FA	inst1579	(r17s_reg[28], pp_reg[572], r18c[26], r18s[27], r18c[27]);
FA	inst1580	(r17s_reg[29], pp_reg[573], r18c[27], r18s[28], r18c[28]);
FA	inst1581	(r17s_reg[30], pp_reg[574], r18c[28], r18s[29], r18c[29]);
FA	inst1582	(rc_last_reg[16], pp_reg[575], r18c[29], r18s[30], r18c[30]);
//Posible pipline
always @(posedge clk) begin
	r18s_reg <= r18s;
	rc_last_reg[17] <= r18c[30];
	ProcConditon_reg[18] <= ProcConditon_reg[17];
end

HA	inst1583	(r18s_reg[1], pp_reg[608], m[19], r19c[0]);
FA	inst1584	(r18s_reg[2], pp_reg[609], r19c[0], r19s[1], r19c[1]);
FA	inst1585	(r18s_reg[3], pp_reg[610], r19c[1], r19s[2], r19c[2]);
FA	inst1586	(r18s_reg[4], pp_reg[611], r19c[2], r19s[3], r19c[3]);
FA	inst1587	(r18s_reg[5], pp_reg[612], r19c[3], r19s[4], r19c[4]);
FA	inst1588	(r18s_reg[6], pp_reg[613], r19c[4], r19s[5], r19c[5]);
FA	inst1589	(r18s_reg[7], pp_reg[614], r19c[5], r19s[6], r19c[6]);
FA	inst1590	(r18s_reg[8], pp_reg[615], r19c[6], r19s[7], r19c[7]);
FA	inst1591	(r18s_reg[9], pp_reg[616], r19c[7], r19s[8], r19c[8]);
FA	inst1592	(r18s_reg[10], pp_reg[617], r19c[8], r19s[9], r19c[9]);
FA	inst1593	(r18s_reg[11], pp_reg[618], r19c[9], r19s[10], r19c[10]);
FA	inst1594	(r18s_reg[12], pp_reg[619], r19c[10], r19s[11], r19c[11]);
FA	inst1595	(r18s_reg[13], pp_reg[620], r19c[11], r19s[12], r19c[12]);
FA	inst1596	(r18s_reg[14], pp_reg[590], r19c[12], r19s[13], r19c[13]);
FA	inst1597	(r18s_reg[15], pp_reg[591], r19c[13], r19s[14], r19c[14]);
FA	inst1598	(r18s_reg[16], pp_reg[592], r19c[14], r19s[15], r19c[15]);
FA	inst1599	(r18s_reg[17], pp_reg[593], r19c[15], r19s[16], r19c[16]);
FA	inst1600	(r18s_reg[18], pp_reg[594], r19c[16], r19s[17], r19c[17]);
FA	inst1601	(r18s_reg[19], pp_reg[595], r19c[17], r19s[18], r19c[18]);
FA	inst1602	(r18s_reg[20], pp_reg[596], r19c[18], r19s[19], r19c[19]);
FA	inst1603	(r18s_reg[21], pp_reg[597], r19c[19], r19s[20], r19c[20]);
FA	inst1604	(r18s_reg[22], pp_reg[598], r19c[20], r19s[21], r19c[21]);
FA	inst1605	(r18s_reg[23], pp_reg[599], r19c[21], r19s[22], r19c[22]);
FA	inst1606	(r18s_reg[24], pp_reg[600], r19c[22], r19s[23], r19c[23]);
FA	inst1607	(r18s_reg[25], pp_reg[601], r19c[23], r19s[24], r19c[24]);
FA	inst1608	(r18s_reg[26], pp_reg[602], r19c[24], r19s[25], r19c[25]);
FA	inst1609	(r18s_reg[27], pp_reg[603], r19c[25], r19s[26], r19c[26]);
FA	inst1610	(r18s_reg[28], pp_reg[604], r19c[26], r19s[27], r19c[27]);
FA	inst1611	(r18s_reg[29], pp_reg[605], r19c[27], r19s[28], r19c[28]);
FA	inst1612	(r18s_reg[30], pp_reg[606], r19c[28], r19s[29], r19c[29]);
FA	inst1613	(rc_last_reg[17], pp_reg[607], r19c[29], r19s[30], r19c[30]);
//Posible pipline
always @(posedge clk) begin
	r19s_reg <= r19s;
	rc_last_reg[18] <= r19c[30];
	ProcConditon_reg[19] <= ProcConditon_reg[18];
end

HA	inst1614	(r19s_reg[1], pp_reg[640], m[20], r20c[0]);
FA	inst1615	(r19s_reg[2], pp_reg[641], r20c[0], r20s[1], r20c[1]);
FA	inst1616	(r19s_reg[3], pp_reg[642], r20c[1], r20s[2], r20c[2]);
FA	inst1617	(r19s_reg[4], pp_reg[643], r20c[2], r20s[3], r20c[3]);
FA	inst1618	(r19s_reg[5], pp_reg[644], r20c[3], r20s[4], r20c[4]);
FA	inst1619	(r19s_reg[6], pp_reg[645], r20c[4], r20s[5], r20c[5]);
FA	inst1620	(r19s_reg[7], pp_reg[646], r20c[5], r20s[6], r20c[6]);
FA	inst1621	(r19s_reg[8], pp_reg[647], r20c[6], r20s[7], r20c[7]);
FA	inst1622	(r19s_reg[9], pp_reg[648], r20c[7], r20s[8], r20c[8]);
FA	inst1623	(r19s_reg[10], pp_reg[649], r20c[8], r20s[9], r20c[9]);
FA	inst1624	(r19s_reg[11], pp_reg[650], r20c[9], r20s[10], r20c[10]);
FA	inst1625	(r19s_reg[12], pp_reg[651], r20c[10], r20s[11], r20c[11]);
FA	inst1626	(r19s_reg[13], pp_reg[621], r20c[11], r20s[12], r20c[12]);
FA	inst1627	(r19s_reg[14], pp_reg[622], r20c[12], r20s[13], r20c[13]);
FA	inst1628	(r19s_reg[15], pp_reg[623], r20c[13], r20s[14], r20c[14]);
FA	inst1629	(r19s_reg[16], pp_reg[624], r20c[14], r20s[15], r20c[15]);
FA	inst1630	(r19s_reg[17], pp_reg[625], r20c[15], r20s[16], r20c[16]);
FA	inst1631	(r19s_reg[18], pp_reg[626], r20c[16], r20s[17], r20c[17]);
FA	inst1632	(r19s_reg[19], pp_reg[627], r20c[17], r20s[18], r20c[18]);
FA	inst1633	(r19s_reg[20], pp_reg[628], r20c[18], r20s[19], r20c[19]);
FA	inst1634	(r19s_reg[21], pp_reg[629], r20c[19], r20s[20], r20c[20]);
FA	inst1635	(r19s_reg[22], pp_reg[630], r20c[20], r20s[21], r20c[21]);
FA	inst1636	(r19s_reg[23], pp_reg[631], r20c[21], r20s[22], r20c[22]);
FA	inst1637	(r19s_reg[24], pp_reg[632], r20c[22], r20s[23], r20c[23]);
FA	inst1638	(r19s_reg[25], pp_reg[633], r20c[23], r20s[24], r20c[24]);
FA	inst1639	(r19s_reg[26], pp_reg[634], r20c[24], r20s[25], r20c[25]);
FA	inst1640	(r19s_reg[27], pp_reg[635], r20c[25], r20s[26], r20c[26]);
FA	inst1641	(r19s_reg[28], pp_reg[636], r20c[26], r20s[27], r20c[27]);
FA	inst1642	(r19s_reg[29], pp_reg[637], r20c[27], r20s[28], r20c[28]);
FA	inst1643	(r19s_reg[30], pp_reg[638], r20c[28], r20s[29], r20c[29]);
FA	inst1644	(rc_last_reg[18], pp_reg[639], r20c[29], r20s[30], r20c[30]);
//Posible pipline
always @(posedge clk) begin
	r20s_reg <= r20s;
	rc_last_reg[19] <= r20c[30];
	ProcConditon_reg[20] <= ProcConditon_reg[19];
end

HA	inst1645	(r20s_reg[1], pp_reg[672], m[21], r21c[0]);
FA	inst1646	(r20s_reg[2], pp_reg[673], r21c[0], r21s[1], r21c[1]);
FA	inst1647	(r20s_reg[3], pp_reg[674], r21c[1], r21s[2], r21c[2]);
FA	inst1648	(r20s_reg[4], pp_reg[675], r21c[2], r21s[3], r21c[3]);
FA	inst1649	(r20s_reg[5], pp_reg[676], r21c[3], r21s[4], r21c[4]);
FA	inst1650	(r20s_reg[6], pp_reg[677], r21c[4], r21s[5], r21c[5]);
FA	inst1651	(r20s_reg[7], pp_reg[678], r21c[5], r21s[6], r21c[6]);
FA	inst1652	(r20s_reg[8], pp_reg[679], r21c[6], r21s[7], r21c[7]);
FA	inst1653	(r20s_reg[9], pp_reg[680], r21c[7], r21s[8], r21c[8]);
FA	inst1654	(r20s_reg[10], pp_reg[681], r21c[8], r21s[9], r21c[9]);
FA	inst1655	(r20s_reg[11], pp_reg[682], r21c[9], r21s[10], r21c[10]);
FA	inst1656	(r20s_reg[12], pp_reg[652], r21c[10], r21s[11], r21c[11]);
FA	inst1657	(r20s_reg[13], pp_reg[653], r21c[11], r21s[12], r21c[12]);
FA	inst1658	(r20s_reg[14], pp_reg[654], r21c[12], r21s[13], r21c[13]);
FA	inst1659	(r20s_reg[15], pp_reg[655], r21c[13], r21s[14], r21c[14]);
FA	inst1660	(r20s_reg[16], pp_reg[656], r21c[14], r21s[15], r21c[15]);
FA	inst1661	(r20s_reg[17], pp_reg[657], r21c[15], r21s[16], r21c[16]);
FA	inst1662	(r20s_reg[18], pp_reg[658], r21c[16], r21s[17], r21c[17]);
FA	inst1663	(r20s_reg[19], pp_reg[659], r21c[17], r21s[18], r21c[18]);
FA	inst1664	(r20s_reg[20], pp_reg[660], r21c[18], r21s[19], r21c[19]);
FA	inst1665	(r20s_reg[21], pp_reg[661], r21c[19], r21s[20], r21c[20]);
FA	inst1666	(r20s_reg[22], pp_reg[662], r21c[20], r21s[21], r21c[21]);
FA	inst1667	(r20s_reg[23], pp_reg[663], r21c[21], r21s[22], r21c[22]);
FA	inst1668	(r20s_reg[24], pp_reg[664], r21c[22], r21s[23], r21c[23]);
FA	inst1669	(r20s_reg[25], pp_reg[665], r21c[23], r21s[24], r21c[24]);
FA	inst1670	(r20s_reg[26], pp_reg[666], r21c[24], r21s[25], r21c[25]);
FA	inst1671	(r20s_reg[27], pp_reg[667], r21c[25], r21s[26], r21c[26]);
FA	inst1672	(r20s_reg[28], pp_reg[668], r21c[26], r21s[27], r21c[27]);
FA	inst1673	(r20s_reg[29], pp_reg[669], r21c[27], r21s[28], r21c[28]);
FA	inst1674	(r20s_reg[30], pp_reg[670], r21c[28], r21s[29], r21c[29]);
FA	inst1675	(rc_last_reg[19], pp_reg[671], r21c[29], r21s[30], r21c[30]);
//Posible pipline
always @(posedge clk) begin
	r21s_reg <= r21s;
	rc_last_reg[20] <= r21c[30];
	ProcConditon_reg[21] <= ProcConditon_reg[20];
end

HA	inst1676	(r21s_reg[1], pp_reg[704], m[22], r22c[0]);
FA	inst1677	(r21s_reg[2], pp_reg[705], r22c[0], r22s[1], r22c[1]);
FA	inst1678	(r21s_reg[3], pp_reg[706], r22c[1], r22s[2], r22c[2]);
FA	inst1679	(r21s_reg[4], pp_reg[707], r22c[2], r22s[3], r22c[3]);
FA	inst1680	(r21s_reg[5], pp_reg[708], r22c[3], r22s[4], r22c[4]);
FA	inst1681	(r21s_reg[6], pp_reg[709], r22c[4], r22s[5], r22c[5]);
FA	inst1682	(r21s_reg[7], pp_reg[710], r22c[5], r22s[6], r22c[6]);
FA	inst1683	(r21s_reg[8], pp_reg[711], r22c[6], r22s[7], r22c[7]);
FA	inst1684	(r21s_reg[9], pp_reg[712], r22c[7], r22s[8], r22c[8]);
FA	inst1685	(r21s_reg[10], pp_reg[713], r22c[8], r22s[9], r22c[9]);
FA	inst1686	(r21s_reg[11], pp_reg[683], r22c[9], r22s[10], r22c[10]);
FA	inst1687	(r21s_reg[12], pp_reg[684], r22c[10], r22s[11], r22c[11]);
FA	inst1688	(r21s_reg[13], pp_reg[685], r22c[11], r22s[12], r22c[12]);
FA	inst1689	(r21s_reg[14], pp_reg[686], r22c[12], r22s[13], r22c[13]);
FA	inst1690	(r21s_reg[15], pp_reg[687], r22c[13], r22s[14], r22c[14]);
FA	inst1691	(r21s_reg[16], pp_reg[688], r22c[14], r22s[15], r22c[15]);
FA	inst1692	(r21s_reg[17], pp_reg[689], r22c[15], r22s[16], r22c[16]);
FA	inst1693	(r21s_reg[18], pp_reg[690], r22c[16], r22s[17], r22c[17]);
FA	inst1694	(r21s_reg[19], pp_reg[691], r22c[17], r22s[18], r22c[18]);
FA	inst1695	(r21s_reg[20], pp_reg[692], r22c[18], r22s[19], r22c[19]);
FA	inst1696	(r21s_reg[21], pp_reg[693], r22c[19], r22s[20], r22c[20]);
FA	inst1697	(r21s_reg[22], pp_reg[694], r22c[20], r22s[21], r22c[21]);
FA	inst1698	(r21s_reg[23], pp_reg[695], r22c[21], r22s[22], r22c[22]);
FA	inst1699	(r21s_reg[24], pp_reg[696], r22c[22], r22s[23], r22c[23]);
FA	inst1700	(r21s_reg[25], pp_reg[697], r22c[23], r22s[24], r22c[24]);
FA	inst1701	(r21s_reg[26], pp_reg[698], r22c[24], r22s[25], r22c[25]);
FA	inst1702	(r21s_reg[27], pp_reg[699], r22c[25], r22s[26], r22c[26]);
FA	inst1703	(r21s_reg[28], pp_reg[700], r22c[26], r22s[27], r22c[27]);
FA	inst1704	(r21s_reg[29], pp_reg[701], r22c[27], r22s[28], r22c[28]);
FA	inst1705	(r21s_reg[30], pp_reg[702], r22c[28], r22s[29], r22c[29]);
FA	inst1706	(rc_last_reg[20], pp_reg[703], r22c[29], r22s[30], r22c[30]);
//Posible pipline
always @(posedge clk) begin
	r22s_reg <= r22s;
	rc_last_reg[21] <= r22c[30];
	ProcConditon_reg[22] <= ProcConditon_reg[20];
end

HA	inst1707	(r22s[1], pp_reg[736], m[23], r23c[0]);
FA	inst1708	(r22s[2], pp_reg[737], r23c[0], r23s[1], r23c[1]);
FA	inst1709	(r22s[3], pp_reg[738], r23c[1], r23s[2], r23c[2]);
FA	inst1710	(r22s[4], pp_reg[739], r23c[2], r23s[3], r23c[3]);
FA	inst1711	(r22s[5], pp_reg[740], r23c[3], r23s[4], r23c[4]);
FA	inst1712	(r22s[6], pp_reg[741], r23c[4], r23s[5], r23c[5]);
FA	inst1713	(r22s[7], pp_reg[742], r23c[5], r23s[6], r23c[6]);
FA	inst1714	(r22s[8], pp_reg[743], r23c[6], r23s[7], r23c[7]);
FA	inst1715	(r22s[9], pp_reg[744], r23c[7], r23s[8], r23c[8]);
FA	inst1716	(r22s[10], pp_reg[714], r23c[8], r23s[9], r23c[9]);
FA	inst1717	(r22s[11], pp_reg[715], r23c[9], r23s[10], r23c[10]);
FA	inst1718	(r22s[12], pp_reg[716], r23c[10], r23s[11], r23c[11]);
FA	inst1719	(r22s[13], pp_reg[717], r23c[11], r23s[12], r23c[12]);
FA	inst1720	(r22s[14], pp_reg[718], r23c[12], r23s[13], r23c[13]);
FA	inst1721	(r22s[15], pp_reg[719], r23c[13], r23s[14], r23c[14]);
FA	inst1722	(r22s[16], pp_reg[720], r23c[14], r23s[15], r23c[15]);
FA	inst1723	(r22s[17], pp_reg[721], r23c[15], r23s[16], r23c[16]);
FA	inst1724	(r22s[18], pp_reg[722], r23c[16], r23s[17], r23c[17]);
FA	inst1725	(r22s[19], pp_reg[723], r23c[17], r23s[18], r23c[18]);
FA	inst1726	(r22s[20], pp_reg[724], r23c[18], r23s[19], r23c[19]);
FA	inst1727	(r22s[21], pp_reg[725], r23c[19], r23s[20], r23c[20]);
FA	inst1728	(r22s[22], pp_reg[726], r23c[20], r23s[21], r23c[21]);
FA	inst1729	(r22s[23], pp_reg[727], r23c[21], r23s[22], r23c[22]);
FA	inst1730	(r22s[24], pp_reg[728], r23c[22], r23s[23], r23c[23]);
FA	inst1731	(r22s[25], pp_reg[729], r23c[23], r23s[24], r23c[24]);
FA	inst1732	(r22s[26], pp_reg[730], r23c[24], r23s[25], r23c[25]);
FA	inst1733	(r22s[27], pp_reg[731], r23c[25], r23s[26], r23c[26]);
FA	inst1734	(r22s[28], pp_reg[732], r23c[26], r23s[27], r23c[27]);
FA	inst1735	(r22s[29], pp_reg[733], r23c[27], r23s[28], r23c[28]);
FA	inst1736	(r22s[30], pp_reg[734], r23c[28], r23s[29], r23c[29]);
FA	inst1737	(r22c[30], pp_reg[735], r23c[29], r23s[30], r23c[30]);
//Posible pipline

always @(posedge clk) begin
	r23s_reg <= r23s;
	rc_last_reg[22] <= r23c[30];
	ProcConditon_reg[23] <= ProcConditon_reg[22];
end

HA	inst1738	(r23s_reg[1], pp_reg[768], m[24], r24c[0]);
FA	inst1739	(r23s_reg[2], pp_reg[769], r24c[0], r24s[1], r24c[1]);
FA	inst1740	(r23s_reg[3], pp_reg[770], r24c[1], r24s[2], r24c[2]);
FA	inst1741	(r23s_reg[4], pp_reg[771], r24c[2], r24s[3], r24c[3]);
FA	inst1742	(r23s_reg[5], pp_reg[772], r24c[3], r24s[4], r24c[4]);
FA	inst1743	(r23s_reg[6], pp_reg[773], r24c[4], r24s[5], r24c[5]);
FA	inst1744	(r23s_reg[7], pp_reg[774], r24c[5], r24s[6], r24c[6]);
FA	inst1745	(r23s_reg[8], pp_reg[775], r24c[6], r24s[7], r24c[7]);
FA	inst1746	(r23s_reg[9], pp_reg[745], r24c[7], r24s[8], r24c[8]);
FA	inst1747	(r23s_reg[10], pp_reg[746], r24c[8], r24s[9], r24c[9]);
FA	inst1748	(r23s_reg[11], pp_reg[747], r24c[9], r24s[10], r24c[10]);
FA	inst1749	(r23s_reg[12], pp_reg[748], r24c[10], r24s[11], r24c[11]);
FA	inst1750	(r23s_reg[13], pp_reg[749], r24c[11], r24s[12], r24c[12]);
FA	inst1751	(r23s_reg[14], pp_reg[750], r24c[12], r24s[13], r24c[13]);
FA	inst1752	(r23s_reg[15], pp_reg[751], r24c[13], r24s[14], r24c[14]);
FA	inst1753	(r23s_reg[16], pp_reg[752], r24c[14], r24s[15], r24c[15]);
FA	inst1754	(r23s_reg[17], pp_reg[753], r24c[15], r24s[16], r24c[16]);
FA	inst1755	(r23s_reg[18], pp_reg[754], r24c[16], r24s[17], r24c[17]);
FA	inst1756	(r23s_reg[19], pp_reg[755], r24c[17], r24s[18], r24c[18]);
FA	inst1757	(r23s_reg[20], pp_reg[756], r24c[18], r24s[19], r24c[19]);
FA	inst1758	(r23s_reg[21], pp_reg[757], r24c[19], r24s[20], r24c[20]);
FA	inst1759	(r23s_reg[22], pp_reg[758], r24c[20], r24s[21], r24c[21]);
FA	inst1760	(r23s_reg[23], pp_reg[759], r24c[21], r24s[22], r24c[22]);
FA	inst1761	(r23s_reg[24], pp_reg[760], r24c[22], r24s[23], r24c[23]);
FA	inst1762	(r23s_reg[25], pp_reg[761], r24c[23], r24s[24], r24c[24]);
FA	inst1763	(r23s_reg[26], pp_reg[762], r24c[24], r24s[25], r24c[25]);
FA	inst1764	(r23s_reg[27], pp_reg[763], r24c[25], r24s[26], r24c[26]);
FA	inst1765	(r23s_reg[28], pp_reg[764], r24c[26], r24s[27], r24c[27]);
FA	inst1766	(r23s_reg[29], pp_reg[765], r24c[27], r24s[28], r24c[28]);
FA	inst1767	(r23s_reg[30], pp_reg[766], r24c[28], r24s[29], r24c[29]);
FA	inst1768	(rc_last_reg[22], pp_reg[767], r24c[29], r24s[30], r24c[30]);
//Posible pipline
always @(posedge clk) begin
	r24s_reg <= r24s;
	rc_last_reg[23] <= r24c[30];
	ProcConditon_reg[24] <= ProcConditon_reg[23];
end

HA	inst1769	(r24s_reg[1], pp_reg[800], m[25], r25c[0]);
FA	inst1770	(r24s_reg[2], pp_reg[801], r25c[0], r25s[1], r25c[1]);
FA	inst1771	(r24s_reg[3], pp_reg[802], r25c[1], r25s[2], r25c[2]);
FA	inst1772	(r24s_reg[4], pp_reg[803], r25c[2], r25s[3], r25c[3]);
FA	inst1773	(r24s_reg[5], pp_reg[804], r25c[3], r25s[4], r25c[4]);
FA	inst1774	(r24s_reg[6], pp_reg[805], r25c[4], r25s[5], r25c[5]);
FA	inst1775	(r24s_reg[7], pp_reg[806], r25c[5], r25s[6], r25c[6]);
FA	inst1776	(r24s_reg[8], pp_reg[776], r25c[6], r25s[7], r25c[7]);
FA	inst1777	(r24s_reg[9], pp_reg[777], r25c[7], r25s[8], r25c[8]);
FA	inst1778	(r24s_reg[10], pp_reg[778], r25c[8], r25s[9], r25c[9]);
FA	inst1779	(r24s_reg[11], pp_reg[779], r25c[9], r25s[10], r25c[10]);
FA	inst1780	(r24s_reg[12], pp_reg[780], r25c[10], r25s[11], r25c[11]);
FA	inst1781	(r24s_reg[13], pp_reg[781], r25c[11], r25s[12], r25c[12]);
FA	inst1782	(r24s_reg[14], pp_reg[782], r25c[12], r25s[13], r25c[13]);
FA	inst1783	(r24s_reg[15], pp_reg[783], r25c[13], r25s[14], r25c[14]);
FA	inst1784	(r24s_reg[16], pp_reg[784], r25c[14], r25s[15], r25c[15]);
FA	inst1785	(r24s_reg[17], pp_reg[785], r25c[15], r25s[16], r25c[16]);
FA	inst1786	(r24s_reg[18], pp_reg[786], r25c[16], r25s[17], r25c[17]);
FA	inst1787	(r24s_reg[19], pp_reg[787], r25c[17], r25s[18], r25c[18]);
FA	inst1788	(r24s_reg[20], pp_reg[788], r25c[18], r25s[19], r25c[19]);
FA	inst1789	(r24s_reg[21], pp_reg[789], r25c[19], r25s[20], r25c[20]);
FA	inst1790	(r24s_reg[22], pp_reg[790], r25c[20], r25s[21], r25c[21]);
FA	inst1791	(r24s_reg[23], pp_reg[791], r25c[21], r25s[22], r25c[22]);
FA	inst1792	(r24s_reg[24], pp_reg[792], r25c[22], r25s[23], r25c[23]);
FA	inst1793	(r24s_reg[25], pp_reg[793], r25c[23], r25s[24], r25c[24]);
FA	inst1794	(r24s_reg[26], pp_reg[794], r25c[24], r25s[25], r25c[25]);
FA	inst1795	(r24s_reg[27], pp_reg[795], r25c[25], r25s[26], r25c[26]);
FA	inst1796	(r24s_reg[28], pp_reg[796], r25c[26], r25s[27], r25c[27]);
FA	inst1797	(r24s_reg[29], pp_reg[797], r25c[27], r25s[28], r25c[28]);
FA	inst1798	(r24s_reg[30], pp_reg[798], r25c[28], r25s[29], r25c[29]);
FA	inst1799	(rc_last_reg[23], pp_reg[799], r25c[29], r25s[30], r25c[30]);
//Posible pipline
always @(posedge clk) begin
	r25s_reg <= r25s;
	rc_last_reg[24] <= r25c[30];
	ProcConditon_reg[25] <= ProcConditon_reg[24];
end

HA	inst1800	(r25s_reg[1], pp_reg[832], m[26], r26c[0]);
FA	inst1801	(r25s_reg[2], pp_reg[833], r26c[0], r26s[1], r26c[1]);
FA	inst1802	(r25s_reg[3], pp_reg[834], r26c[1], r26s[2], r26c[2]);
FA	inst1803	(r25s_reg[4], pp_reg[835], r26c[2], r26s[3], r26c[3]);
FA	inst1804	(r25s_reg[5], pp_reg[836], r26c[3], r26s[4], r26c[4]);
FA	inst1805	(r25s_reg[6], pp_reg[837], r26c[4], r26s[5], r26c[5]);
FA	inst1806	(r25s_reg[7], pp_reg[807], r26c[5], r26s[6], r26c[6]);
FA	inst1807	(r25s_reg[8], pp_reg[808], r26c[6], r26s[7], r26c[7]);
FA	inst1808	(r25s_reg[9], pp_reg[809], r26c[7], r26s[8], r26c[8]);
FA	inst1809	(r25s_reg[10], pp_reg[810], r26c[8], r26s[9], r26c[9]);
FA	inst1810	(r25s_reg[11], pp_reg[811], r26c[9], r26s[10], r26c[10]);
FA	inst1811	(r25s_reg[12], pp_reg[812], r26c[10], r26s[11], r26c[11]);
FA	inst1812	(r25s_reg[13], pp_reg[813], r26c[11], r26s[12], r26c[12]);
FA	inst1813	(r25s_reg[14], pp_reg[814], r26c[12], r26s[13], r26c[13]);
FA	inst1814	(r25s_reg[15], pp_reg[815], r26c[13], r26s[14], r26c[14]);
FA	inst1815	(r25s_reg[16], pp_reg[816], r26c[14], r26s[15], r26c[15]);
FA	inst1816	(r25s_reg[17], pp_reg[817], r26c[15], r26s[16], r26c[16]);
FA	inst1817	(r25s_reg[18], pp_reg[818], r26c[16], r26s[17], r26c[17]);
FA	inst1818	(r25s_reg[19], pp_reg[819], r26c[17], r26s[18], r26c[18]);
FA	inst1819	(r25s_reg[20], pp_reg[820], r26c[18], r26s[19], r26c[19]);
FA	inst1820	(r25s_reg[21], pp_reg[821], r26c[19], r26s[20], r26c[20]);
FA	inst1821	(r25s_reg[22], pp_reg[822], r26c[20], r26s[21], r26c[21]);
FA	inst1822	(r25s_reg[23], pp_reg[823], r26c[21], r26s[22], r26c[22]);
FA	inst1823	(r25s_reg[24], pp_reg[824], r26c[22], r26s[23], r26c[23]);
FA	inst1824	(r25s_reg[25], pp_reg[825], r26c[23], r26s[24], r26c[24]);
FA	inst1825	(r25s_reg[26], pp_reg[826], r26c[24], r26s[25], r26c[25]);
FA	inst1826	(r25s_reg[27], pp_reg[827], r26c[25], r26s[26], r26c[26]);
FA	inst1827	(r25s_reg[28], pp_reg[828], r26c[26], r26s[27], r26c[27]);
FA	inst1828	(r25s_reg[29], pp_reg[829], r26c[27], r26s[28], r26c[28]);
FA	inst1829	(r25s_reg[30], pp_reg[830], r26c[28], r26s[29], r26c[29]);
FA	inst1830	(rc_last_reg[24], pp_reg[831], r26c[29], r26s[30], r26c[30]);
//Posible pipline
always @(posedge clk) begin
	r26s_reg <= r26s;
	rc_last_reg[25] <= r26c[30];
	ProcConditon_reg[26] <= ProcConditon_reg[25];
end

HA	inst1831	(r26s_reg[1], pp_reg[864], m[27], r27c[0]);
FA	inst1832	(r26s_reg[2], pp_reg[865], r27c[0], r27s[1], r27c[1]);
FA	inst1833	(r26s_reg[3], pp_reg[866], r27c[1], r27s[2], r27c[2]);
FA	inst1834	(r26s_reg[4], pp_reg[867], r27c[2], r27s[3], r27c[3]);
FA	inst1835	(r26s_reg[5], pp_reg[868], r27c[3], r27s[4], r27c[4]);
FA	inst1836	(r26s_reg[6], pp_reg[838], r27c[4], r27s[5], r27c[5]);
FA	inst1837	(r26s_reg[7], pp_reg[839], r27c[5], r27s[6], r27c[6]);
FA	inst1838	(r26s_reg[8], pp_reg[840], r27c[6], r27s[7], r27c[7]);
FA	inst1839	(r26s_reg[9], pp_reg[841], r27c[7], r27s[8], r27c[8]);
FA	inst1840	(r26s_reg[10], pp_reg[842], r27c[8], r27s[9], r27c[9]);
FA	inst1841	(r26s_reg[11], pp_reg[843], r27c[9], r27s[10], r27c[10]);
FA	inst1842	(r26s_reg[12], pp_reg[844], r27c[10], r27s[11], r27c[11]);
FA	inst1843	(r26s_reg[13], pp_reg[845], r27c[11], r27s[12], r27c[12]);
FA	inst1844	(r26s_reg[14], pp_reg[846], r27c[12], r27s[13], r27c[13]);
FA	inst1845	(r26s_reg[15], pp_reg[847], r27c[13], r27s[14], r27c[14]);
FA	inst1846	(r26s_reg[16], pp_reg[848], r27c[14], r27s[15], r27c[15]);
FA	inst1847	(r26s_reg[17], pp_reg[849], r27c[15], r27s[16], r27c[16]);
FA	inst1848	(r26s_reg[18], pp_reg[850], r27c[16], r27s[17], r27c[17]);
FA	inst1849	(r26s_reg[19], pp_reg[851], r27c[17], r27s[18], r27c[18]);
FA	inst1850	(r26s_reg[20], pp_reg[852], r27c[18], r27s[19], r27c[19]);
FA	inst1851	(r26s_reg[21], pp_reg[853], r27c[19], r27s[20], r27c[20]);
FA	inst1852	(r26s_reg[22], pp_reg[854], r27c[20], r27s[21], r27c[21]);
FA	inst1853	(r26s_reg[23], pp_reg[855], r27c[21], r27s[22], r27c[22]);
FA	inst1854	(r26s_reg[24], pp_reg[856], r27c[22], r27s[23], r27c[23]);
FA	inst1855	(r26s_reg[25], pp_reg[857], r27c[23], r27s[24], r27c[24]);
FA	inst1856	(r26s_reg[26], pp_reg[858], r27c[24], r27s[25], r27c[25]);
FA	inst1857	(r26s_reg[27], pp_reg[859], r27c[25], r27s[26], r27c[26]);
FA	inst1858	(r26s_reg[28], pp_reg[860], r27c[26], r27s[27], r27c[27]);
FA	inst1859	(r26s_reg[29], pp_reg[861], r27c[27], r27s[28], r27c[28]);
FA	inst1860	(r26s_reg[30], pp_reg[862], r27c[28], r27s[29], r27c[29]);
FA	inst1861	(rc_last_reg[25], pp_reg[863], r27c[29], r27s[30], r27c[30]);
//Posible pipline
always @(posedge clk) begin
	r27s_reg <= r27s;
	rc_last_reg[26] <= r27c[30];
	ProcConditon_reg[27] <= ProcConditon_reg[26];
end

HA	inst1862	(r27s_reg[1], pp_reg[896], m[28], r28c[0]);
FA	inst1863	(r27s_reg[2], pp_reg[897], r28c[0], r28s[1], r28c[1]);
FA	inst1864	(r27s_reg[3], pp_reg[898], r28c[1], r28s[2], r28c[2]);
FA	inst1865	(r27s_reg[4], pp_reg[899], r28c[2], r28s[3], r28c[3]);
FA	inst1866	(r27s_reg[5], pp_reg[869], r28c[3], r28s[4], r28c[4]);
FA	inst1867	(r27s_reg[6], pp_reg[870], r28c[4], r28s[5], r28c[5]);
FA	inst1868	(r27s_reg[7], pp_reg[871], r28c[5], r28s[6], r28c[6]);
FA	inst1869	(r27s_reg[8], pp_reg[872], r28c[6], r28s[7], r28c[7]);
FA	inst1870	(r27s_reg[9], pp_reg[873], r28c[7], r28s[8], r28c[8]);
FA	inst1871	(r27s_reg[10], pp_reg[874], r28c[8], r28s[9], r28c[9]);
FA	inst1872	(r27s_reg[11], pp_reg[875], r28c[9], r28s[10], r28c[10]);
FA	inst1873	(r27s_reg[12], pp_reg[876], r28c[10], r28s[11], r28c[11]);
FA	inst1874	(r27s_reg[13], pp_reg[877], r28c[11], r28s[12], r28c[12]);
FA	inst1875	(r27s_reg[14], pp_reg[878], r28c[12], r28s[13], r28c[13]);
FA	inst1876	(r27s_reg[15], pp_reg[879], r28c[13], r28s[14], r28c[14]);
FA	inst1877	(r27s_reg[16], pp_reg[880], r28c[14], r28s[15], r28c[15]);
FA	inst1878	(r27s_reg[17], pp_reg[881], r28c[15], r28s[16], r28c[16]);
FA	inst1879	(r27s_reg[18], pp_reg[882], r28c[16], r28s[17], r28c[17]);
FA	inst1880	(r27s_reg[19], pp_reg[883], r28c[17], r28s[18], r28c[18]);
FA	inst1881	(r27s_reg[20], pp_reg[884], r28c[18], r28s[19], r28c[19]);
FA	inst1882	(r27s_reg[21], pp_reg[885], r28c[19], r28s[20], r28c[20]);
FA	inst1883	(r27s_reg[22], pp_reg[886], r28c[20], r28s[21], r28c[21]);
FA	inst1884	(r27s_reg[23], pp_reg[887], r28c[21], r28s[22], r28c[22]);
FA	inst1885	(r27s_reg[24], pp_reg[888], r28c[22], r28s[23], r28c[23]);
FA	inst1886	(r27s_reg[25], pp_reg[889], r28c[23], r28s[24], r28c[24]);
FA	inst1887	(r27s_reg[26], pp_reg[890], r28c[24], r28s[25], r28c[25]);
FA	inst1888	(r27s_reg[27], pp_reg[891], r28c[25], r28s[26], r28c[26]);
FA	inst1889	(r27s_reg[28], pp_reg[892], r28c[26], r28s[27], r28c[27]);
FA	inst1890	(r27s_reg[29], pp_reg[893], r28c[27], r28s[28], r28c[28]);
FA	inst1891	(r27s_reg[30], pp_reg[894], r28c[28], r28s[29], r28c[29]);
FA	inst1892	(rc_last_reg[26], pp_reg[895], r28c[29], r28s[30], r28c[30]);
//Posible pipline
always @(posedge clk) begin
	r28s_reg <= r28s;
	rc_last_reg[27] <= r28c[30];
	ProcConditon_reg[28] <= ProcConditon_reg[27];
end

HA	inst1893	(r28s_reg[1], pp_reg[928], m[29], r29c[0]);
FA	inst1894	(r28s_reg[2], pp_reg[929], r29c[0], r29s[1], r29c[1]);
FA	inst1895	(r28s_reg[3], pp_reg[930], r29c[1], r29s[2], r29c[2]);
FA	inst1896	(r28s_reg[4], pp_reg[900], r29c[2], r29s[3], r29c[3]);
FA	inst1897	(r28s_reg[5], pp_reg[901], r29c[3], r29s[4], r29c[4]);
FA	inst1898	(r28s_reg[6], pp_reg[902], r29c[4], r29s[5], r29c[5]);
FA	inst1899	(r28s_reg[7], pp_reg[903], r29c[5], r29s[6], r29c[6]);
FA	inst1900	(r28s_reg[8], pp_reg[904], r29c[6], r29s[7], r29c[7]);
FA	inst1901	(r28s_reg[9], pp_reg[905], r29c[7], r29s[8], r29c[8]);
FA	inst1902	(r28s_reg[10], pp_reg[906], r29c[8], r29s[9], r29c[9]);
FA	inst1903	(r28s_reg[11], pp_reg[907], r29c[9], r29s[10], r29c[10]);
FA	inst1904	(r28s_reg[12], pp_reg[908], r29c[10], r29s[11], r29c[11]);
FA	inst1905	(r28s_reg[13], pp_reg[909], r29c[11], r29s[12], r29c[12]);
FA	inst1906	(r28s_reg[14], pp_reg[910], r29c[12], r29s[13], r29c[13]);
FA	inst1907	(r28s_reg[15], pp_reg[911], r29c[13], r29s[14], r29c[14]);
FA	inst1908	(r28s_reg[16], pp_reg[912], r29c[14], r29s[15], r29c[15]);
FA	inst1909	(r28s_reg[17], pp_reg[913], r29c[15], r29s[16], r29c[16]);
FA	inst1910	(r28s_reg[18], pp_reg[914], r29c[16], r29s[17], r29c[17]);
FA	inst1911	(r28s_reg[19], pp_reg[915], r29c[17], r29s[18], r29c[18]);
FA	inst1912	(r28s_reg[20], pp_reg[916], r29c[18], r29s[19], r29c[19]);
FA	inst1913	(r28s_reg[21], pp_reg[917], r29c[19], r29s[20], r29c[20]);
FA	inst1914	(r28s_reg[22], pp_reg[918], r29c[20], r29s[21], r29c[21]);
FA	inst1915	(r28s_reg[23], pp_reg[919], r29c[21], r29s[22], r29c[22]);
FA	inst1916	(r28s_reg[24], pp_reg[920], r29c[22], r29s[23], r29c[23]);
FA	inst1917	(r28s_reg[25], pp_reg[921], r29c[23], r29s[24], r29c[24]);
FA	inst1918	(r28s_reg[26], pp_reg[922], r29c[24], r29s[25], r29c[25]);
FA	inst1919	(r28s_reg[27], pp_reg[923], r29c[25], r29s[26], r29c[26]);
FA	inst1920	(r28s_reg[28], pp_reg[924], r29c[26], r29s[27], r29c[27]);
FA	inst1921	(r28s_reg[29], pp_reg[925], r29c[27], r29s[28], r29c[28]);
FA	inst1922	(r28s_reg[30], pp_reg[926], r29c[28], r29s[29], r29c[29]);
FA	inst1923	(rc_last_reg[27], pp_reg[927], r29c[29], r29s[30], r29c[30]);
//Posible pipline
always @(posedge clk) begin
	r29s_reg <= r29s;
	rc_last_reg[28] <= r29c[30];
	ProcConditon_reg[29] <= ProcConditon_reg[28];
end


HA	inst1924	(r29s_reg[1], pp_reg[960], m[30], r30c[0]);
FA	inst1925	(r29s_reg[2], pp_reg[961], r30c[0], r30s[1], r30c[1]);
FA	inst1926	(r29s_reg[3], pp_reg[931], r30c[1], r30s[2], r30c[2]);
FA	inst1927	(r29s_reg[4], pp_reg[932], r30c[2], r30s[3], r30c[3]);
FA	inst1928	(r29s_reg[5], pp_reg[933], r30c[3], r30s[4], r30c[4]);
FA	inst1929	(r29s_reg[6], pp_reg[934], r30c[4], r30s[5], r30c[5]);
FA	inst1930	(r29s_reg[7], pp_reg[935], r30c[5], r30s[6], r30c[6]);
FA	inst1931	(r29s_reg[8], pp_reg[936], r30c[6], r30s[7], r30c[7]);
FA	inst1932	(r29s_reg[9], pp_reg[937], r30c[7], r30s[8], r30c[8]);
FA	inst1933	(r29s_reg[10], pp_reg[938], r30c[8], r30s[9], r30c[9]);
FA	inst1934	(r29s_reg[11], pp_reg[939], r30c[9], r30s[10], r30c[10]);
FA	inst1935	(r29s_reg[12], pp_reg[940], r30c[10], r30s[11], r30c[11]);
FA	inst1936	(r29s_reg[13], pp_reg[941], r30c[11], r30s[12], r30c[12]);
FA	inst1937	(r29s_reg[14], pp_reg[942], r30c[12], r30s[13], r30c[13]);
FA	inst1938	(r29s_reg[15], pp_reg[943], r30c[13], r30s[14], r30c[14]);
FA	inst1939	(r29s_reg[16], pp_reg[944], r30c[14], r30s[15], r30c[15]);
FA	inst1940	(r29s_reg[17], pp_reg[945], r30c[15], r30s[16], r30c[16]);
FA	inst1941	(r29s_reg[18], pp_reg[946], r30c[16], r30s[17], r30c[17]);
FA	inst1942	(r29s_reg[19], pp_reg[947], r30c[17], r30s[18], r30c[18]);
FA	inst1943	(r29s_reg[20], pp_reg[948], r30c[18], r30s[19], r30c[19]);
FA	inst1944	(r29s_reg[21], pp_reg[949], r30c[19], r30s[20], r30c[20]);
FA	inst1945	(r29s_reg[22], pp_reg[950], r30c[20], r30s[21], r30c[21]);
FA	inst1946	(r29s_reg[23], pp_reg[951], r30c[21], r30s[22], r30c[22]);
FA	inst1947	(r29s_reg[24], pp_reg[952], r30c[22], r30s[23], r30c[23]);
FA	inst1948	(r29s_reg[25], pp_reg[953], r30c[23], r30s[24], r30c[24]);
FA	inst1949	(r29s_reg[26], pp_reg[954], r30c[24], r30s[25], r30c[25]);
FA	inst1950	(r29s_reg[27], pp_reg[955], r30c[25], r30s[26], r30c[26]);
FA	inst1951	(r29s_reg[28], pp_reg[956], r30c[26], r30s[27], r30c[27]);
FA	inst1952	(r29s_reg[29], pp_reg[957], r30c[27], r30s[28], r30c[28]);
FA	inst1953	(r29s_reg[30], pp_reg[958], r30c[28], r30s[29], r30c[29]);
FA	inst1954	(rc_last_reg[28], pp_reg[959], r30c[29], r30s[30], r30c[30]);
//Posible pipline
always @(posedge clk) begin
	r30s_reg <= r30s;
	rc_last_reg[29] <= r30c[30];
	ProcConditon_reg[30] <= ProcConditon_reg[29];
end

HA	inst1955	(r30s_reg[1], pp_reg[992], m[31], r31c[0]);
FA	inst1956	(r30s_reg[2], pp_reg[962], r31c[0], r31s[1], r31c[1]);
FA	inst1957	(r30s_reg[3], pp_reg[963], r31c[1], r31s[2], r31c[2]);
FA	inst1958	(r30s_reg[4], pp_reg[964], r31c[2], r31s[3], r31c[3]);
FA	inst1959	(r30s_reg[5], pp_reg[965], r31c[3], r31s[4], r31c[4]);
FA	inst1960	(r30s_reg[6], pp_reg[966], r31c[4], r31s[5], r31c[5]);
FA	inst1961	(r30s_reg[7], pp_reg[967], r31c[5], r31s[6], r31c[6]);
FA	inst1962	(r30s_reg[8], pp_reg[968], r31c[6], r31s[7], r31c[7]);
FA	inst1963	(r30s_reg[9], pp_reg[969], r31c[7], r31s[8], r31c[8]);
FA	inst1964	(r30s_reg[10], pp_reg[970], r31c[8], r31s[9], r31c[9]);
FA	inst1965	(r30s_reg[11], pp_reg[971], r31c[9], r31s[10], r31c[10]);
FA	inst1966	(r30s_reg[12], pp_reg[972], r31c[10], r31s[11], r31c[11]);
FA	inst1967	(r30s_reg[13], pp_reg[973], r31c[11], r31s[12], r31c[12]);
FA	inst1968	(r30s_reg[14], pp_reg[974], r31c[12], r31s[13], r31c[13]);
FA	inst1969	(r30s_reg[15], pp_reg[975], r31c[13], r31s[14], r31c[14]);
FA	inst1970	(r30s_reg[16], pp_reg[976], r31c[14], r31s[15], r31c[15]);
FA	inst1971	(r30s_reg[17], pp_reg[977], r31c[15], r31s[16], r31c[16]);
FA	inst1972	(r30s_reg[18], pp_reg[978], r31c[16], r31s[17], r31c[17]);
FA	inst1973	(r30s_reg[19], pp_reg[979], r31c[17], r31s[18], r31c[18]);
FA	inst1974	(r30s_reg[20], pp_reg[980], r31c[18], r31s[19], r31c[19]);
FA	inst1975	(r30s_reg[21], pp_reg[981], r31c[19], r31s[20], r31c[20]);
FA	inst1976	(r30s_reg[22], pp_reg[982], r31c[20], r31s[21], r31c[21]);
FA	inst1977	(r30s_reg[23], pp_reg[983], r31c[21], r31s[22], r31c[22]);
FA	inst1978	(r30s_reg[24], pp_reg[984], r31c[22], r31s[23], r31c[23]);
FA	inst1979	(r30s_reg[25], pp_reg[985], r31c[23], r31s[24], r31c[24]);
FA	inst1980	(r30s_reg[26], pp_reg[986], r31c[24], r31s[25], r31c[25]);
FA	inst1981	(r30s_reg[27], pp_reg[987], r31c[25], r31s[26], r31c[26]);
FA	inst1982	(r30s_reg[28], pp_reg[988], r31c[26], r31s[27], r31c[27]);
FA	inst1983	(r30s_reg[29], pp_reg[989], r31c[27], r31s[28], r31c[28]);
FA	inst1984	(r30s_reg[30], pp_reg[990], r31c[28], r31s[29], r31c[29]);
FA	inst1985	(rc_last_reg[29], pp_reg[991], r31c[29], r31s[30], r31c[30]);
//Posible pipline
always @(posedge clk) begin
	r31s_reg <= r31s;
	rc_last_reg[30] <= r31c[30];
	PDone_out <= ProcConditon_reg[30];
end

HA	inst1986	(r31s_reg[1], pp_reg[993], m[32], r32c[0]);
FA	inst1987	(r31s_reg[2], pp_reg[994], r32c[0], m[33], r32c[1]);
FA	inst1988	(r31s_reg[3], pp_reg[995], r32c[1], m[34], r32c[2]);
FA	inst1989	(r31s_reg[4], pp_reg[996], r32c[2], m[35], r32c[3]);
FA	inst1990	(r31s_reg[5], pp_reg[997], r32c[3], m[36], r32c[4]);
FA	inst1991	(r31s_reg[6], pp_reg[998], r32c[4], m[37], r32c[5]);
FA	inst1992	(r31s_reg[7], pp_reg[999], r32c[5], m[38], r32c[6]);
FA	inst1993	(r31s_reg[8], pp_reg[1000], r32c[6], m[39], r32c[7]);
FA	inst1994	(r31s_reg[9], pp_reg[1001], r32c[7], m[40], r32c[8]);
FA	inst1995	(r31s_reg[10], pp_reg[1002], r32c[8], m[41], r32c[9]);
FA	inst1996	(r31s_reg[11], pp_reg[1003], r32c[9], m[42], r32c[10]);
FA	inst1997	(r31s_reg[12], pp_reg[1004], r32c[10], m[43], r32c[11]);
FA	inst1998	(r31s_reg[13], pp_reg[1005], r32c[11], m[44], r32c[12]);
FA	inst1999	(r31s_reg[14], pp_reg[1006], r32c[12], m[45], r32c[13]);
FA	inst2000	(r31s_reg[15], pp_reg[1007], r32c[13], m[46], r32c[14]);
FA	inst2001	(r31s_reg[16], pp_reg[1008], r32c[14], m[47], r32c[15]);
FA	inst2002	(r31s_reg[17], pp_reg[1009], r32c[15], m[48], r32c[16]);
FA	inst2003	(r31s_reg[18], pp_reg[1010], r32c[16], m[49], r32c[17]);
FA	inst2004	(r31s_reg[19], pp_reg[1011], r32c[17], m[50], r32c[18]);
FA	inst2005	(r31s_reg[20], pp_reg[1012], r32c[18], m[51], r32c[19]);
FA	inst2006	(r31s_reg[21], pp_reg[1013], r32c[19], m[52], r32c[20]);
FA	inst2007	(r31s_reg[22], pp_reg[1014], r32c[20], m[53], r32c[21]);
FA	inst2008	(r31s_reg[23], pp_reg[1015], r32c[21], m[54], r32c[22]);
FA	inst2009	(r31s_reg[24], pp_reg[1016], r32c[22], m[55], r32c[23]);
FA	inst2010	(r31s_reg[25], pp_reg[1017], r32c[23], m[56], r32c[24]);
FA	inst2011	(r31s_reg[26], pp_reg[1018], r32c[24], m[57], r32c[25]);
FA	inst2012	(r31s_reg[27], pp_reg[1019], r32c[25], m[58], r32c[26]);
FA	inst2013	(r31s_reg[28], pp_reg[1020], r32c[26], m[59], r32c[27]);
FA	inst2014	(r31s_reg[29], pp_reg[1021], r32c[27], m[60], r32c[28]);
FA	inst2015	(r31s_reg[30], pp_reg[1022], r32c[28], m[61], r32c[29]);
FA	inst2016	(rc_last_reg[30], pp_reg[1023], r32c[29], m[62], m[63]);
endmodule
